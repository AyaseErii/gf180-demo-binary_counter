magic
tech gf180mcuC
magscale 1 10
timestamp 1669906326
<< metal1 >>
rect 29026 56590 29038 56642
rect 29090 56639 29102 56642
rect 29922 56639 29934 56642
rect 29090 56593 29934 56639
rect 29090 56590 29102 56593
rect 29922 56590 29934 56593
rect 29986 56590 29998 56642
rect 52322 56590 52334 56642
rect 52386 56639 52398 56642
rect 52994 56639 53006 56642
rect 52386 56593 53006 56639
rect 52386 56590 52398 56593
rect 52994 56590 53006 56593
rect 53058 56590 53070 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 8318 56306 8370 56318
rect 8318 56242 8370 56254
rect 19294 56306 19346 56318
rect 19294 56242 19346 56254
rect 31390 56306 31442 56318
rect 31390 56242 31442 56254
rect 34750 56306 34802 56318
rect 34750 56242 34802 56254
rect 37438 56306 37490 56318
rect 37438 56242 37490 56254
rect 46174 56306 46226 56318
rect 46174 56242 46226 56254
rect 52110 56306 52162 56318
rect 52110 56242 52162 56254
rect 55134 56306 55186 56318
rect 55134 56242 55186 56254
rect 19742 56194 19794 56206
rect 2594 56142 2606 56194
rect 2658 56142 2670 56194
rect 6066 56142 6078 56194
rect 6130 56142 6142 56194
rect 11330 56142 11342 56194
rect 11394 56142 11406 56194
rect 19742 56130 19794 56142
rect 20078 56194 20130 56206
rect 31838 56194 31890 56206
rect 23426 56142 23438 56194
rect 23490 56142 23502 56194
rect 26114 56142 26126 56194
rect 26178 56142 26190 56194
rect 20078 56130 20130 56142
rect 31838 56130 31890 56142
rect 35198 56194 35250 56206
rect 35198 56130 35250 56142
rect 35534 56194 35586 56206
rect 35534 56130 35586 56142
rect 37886 56194 37938 56206
rect 37886 56130 37938 56142
rect 38222 56194 38274 56206
rect 46622 56194 46674 56206
rect 42130 56142 42142 56194
rect 42194 56142 42206 56194
rect 38222 56130 38274 56142
rect 46622 56130 46674 56142
rect 52782 56194 52834 56206
rect 52782 56130 52834 56142
rect 55582 56194 55634 56206
rect 55582 56130 55634 56142
rect 55918 56194 55970 56206
rect 57698 56142 57710 56194
rect 57762 56142 57774 56194
rect 55918 56130 55970 56142
rect 7534 56082 7586 56094
rect 25342 56082 25394 56094
rect 49534 56082 49586 56094
rect 3490 56030 3502 56082
rect 3554 56030 3566 56082
rect 6962 56030 6974 56082
rect 7026 56030 7038 56082
rect 12226 56030 12238 56082
rect 12290 56030 12302 56082
rect 18722 56030 18734 56082
rect 18786 56030 18798 56082
rect 24098 56030 24110 56082
rect 24162 56030 24174 56082
rect 26786 56030 26798 56082
rect 26850 56030 26862 56082
rect 29250 56030 29262 56082
rect 29314 56030 29326 56082
rect 32050 56030 32062 56082
rect 32114 56030 32126 56082
rect 41234 56030 41246 56082
rect 41298 56030 41310 56082
rect 46834 56030 46846 56082
rect 46898 56030 46910 56082
rect 49970 56030 49982 56082
rect 50034 56030 50046 56082
rect 52994 56030 53006 56082
rect 53058 56030 53070 56082
rect 56802 56030 56814 56082
rect 56866 56030 56878 56082
rect 7534 56018 7586 56030
rect 25342 56018 25394 56030
rect 49534 56018 49586 56030
rect 4062 55970 4114 55982
rect 4062 55906 4114 55918
rect 12798 55970 12850 55982
rect 20638 55970 20690 55982
rect 17714 55918 17726 55970
rect 17778 55918 17790 55970
rect 12798 55906 12850 55918
rect 20638 55906 20690 55918
rect 22654 55970 22706 55982
rect 22654 55906 22706 55918
rect 28590 55970 28642 55982
rect 40350 55970 40402 55982
rect 29922 55918 29934 55970
rect 29986 55918 29998 55970
rect 50642 55918 50654 55970
rect 50706 55918 50718 55970
rect 28590 55906 28642 55918
rect 40350 55906 40402 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 55794 55470 55806 55522
rect 55858 55519 55870 55522
rect 56578 55519 56590 55522
rect 55858 55473 56590 55519
rect 55858 55470 55870 55473
rect 56578 55470 56590 55473
rect 56642 55470 56654 55522
rect 57810 55358 57822 55410
rect 57874 55358 57886 55410
rect 11342 55298 11394 55310
rect 10770 55246 10782 55298
rect 10834 55246 10846 55298
rect 11342 55234 11394 55246
rect 15822 55298 15874 55310
rect 16258 55246 16270 55298
rect 16322 55246 16334 55298
rect 56802 55246 56814 55298
rect 56866 55246 56878 55298
rect 15822 55234 15874 55246
rect 1822 55186 1874 55198
rect 1822 55122 1874 55134
rect 2158 55074 2210 55086
rect 2158 55010 2210 55022
rect 7646 55074 7698 55086
rect 11902 55074 11954 55086
rect 8306 55022 8318 55074
rect 8370 55022 8382 55074
rect 7646 55010 7698 55022
rect 11902 55010 11954 55022
rect 12350 55074 12402 55086
rect 19294 55074 19346 55086
rect 18722 55022 18734 55074
rect 18786 55022 18798 55074
rect 12350 55010 12402 55022
rect 19294 55010 19346 55022
rect 19854 55074 19906 55086
rect 19854 55010 19906 55022
rect 20302 55074 20354 55086
rect 20302 55010 20354 55022
rect 20862 55074 20914 55086
rect 20862 55010 20914 55022
rect 55806 55074 55858 55086
rect 55806 55010 55858 55022
rect 56254 55074 56306 55086
rect 56254 55010 56306 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 1822 54738 1874 54750
rect 58046 54738 58098 54750
rect 23202 54686 23214 54738
rect 23266 54686 23278 54738
rect 1822 54674 1874 54686
rect 58046 54674 58098 54686
rect 20078 54514 20130 54526
rect 20738 54462 20750 54514
rect 20802 54462 20814 54514
rect 20078 54450 20130 54462
rect 11454 54402 11506 54414
rect 11454 54338 11506 54350
rect 12350 54402 12402 54414
rect 12350 54338 12402 54350
rect 19630 54402 19682 54414
rect 19630 54338 19682 54350
rect 24222 54402 24274 54414
rect 24222 54338 24274 54350
rect 27806 54402 27858 54414
rect 27806 54338 27858 54350
rect 29150 54402 29202 54414
rect 29150 54338 29202 54350
rect 30718 54402 30770 54414
rect 30718 54338 30770 54350
rect 23774 54290 23826 54302
rect 23774 54226 23826 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 30270 53954 30322 53966
rect 30270 53890 30322 53902
rect 38894 53954 38946 53966
rect 38894 53890 38946 53902
rect 39790 53954 39842 53966
rect 39790 53890 39842 53902
rect 3726 53842 3778 53854
rect 3726 53778 3778 53790
rect 27470 53842 27522 53854
rect 42366 53842 42418 53854
rect 39218 53790 39230 53842
rect 39282 53790 39294 53842
rect 27470 53778 27522 53790
rect 42366 53778 42418 53790
rect 4622 53730 4674 53742
rect 4050 53678 4062 53730
rect 4114 53678 4126 53730
rect 4622 53666 4674 53678
rect 8654 53730 8706 53742
rect 14478 53730 14530 53742
rect 18734 53730 18786 53742
rect 9090 53678 9102 53730
rect 9154 53678 9166 53730
rect 14802 53678 14814 53730
rect 14866 53678 14878 53730
rect 8654 53666 8706 53678
rect 14478 53666 14530 53678
rect 18734 53666 18786 53678
rect 28702 53730 28754 53742
rect 28702 53666 28754 53678
rect 32510 53730 32562 53742
rect 32510 53666 32562 53678
rect 32622 53730 32674 53742
rect 32622 53666 32674 53678
rect 33070 53730 33122 53742
rect 33070 53666 33122 53678
rect 38446 53730 38498 53742
rect 38446 53666 38498 53678
rect 41582 53730 41634 53742
rect 41582 53666 41634 53678
rect 41918 53730 41970 53742
rect 41918 53666 41970 53678
rect 42142 53730 42194 53742
rect 42142 53666 42194 53678
rect 1822 53618 1874 53630
rect 1822 53554 1874 53566
rect 12126 53618 12178 53630
rect 12126 53554 12178 53566
rect 27358 53618 27410 53630
rect 27358 53554 27410 53566
rect 28814 53618 28866 53630
rect 28814 53554 28866 53566
rect 30382 53618 30434 53630
rect 30382 53554 30434 53566
rect 31054 53618 31106 53630
rect 31054 53554 31106 53566
rect 42814 53618 42866 53630
rect 42814 53554 42866 53566
rect 45614 53618 45666 53630
rect 45614 53554 45666 53566
rect 2158 53506 2210 53518
rect 2158 53442 2210 53454
rect 3838 53506 3890 53518
rect 12686 53506 12738 53518
rect 11554 53454 11566 53506
rect 11618 53454 11630 53506
rect 3838 53442 3890 53454
rect 12686 53442 12738 53454
rect 13806 53506 13858 53518
rect 17950 53506 18002 53518
rect 17378 53454 17390 53506
rect 17442 53454 17454 53506
rect 13806 53442 13858 53454
rect 17950 53442 18002 53454
rect 18286 53506 18338 53518
rect 18286 53442 18338 53454
rect 28254 53506 28306 53518
rect 28254 53442 28306 53454
rect 29486 53506 29538 53518
rect 29486 53442 29538 53454
rect 30942 53506 30994 53518
rect 30942 53442 30994 53454
rect 31502 53506 31554 53518
rect 31502 53442 31554 53454
rect 39118 53506 39170 53518
rect 39118 53442 39170 53454
rect 39902 53506 39954 53518
rect 39902 53442 39954 53454
rect 40014 53506 40066 53518
rect 40014 53442 40066 53454
rect 40686 53506 40738 53518
rect 40686 53442 40738 53454
rect 41470 53506 41522 53518
rect 41470 53442 41522 53454
rect 41694 53506 41746 53518
rect 41694 53442 41746 53454
rect 45502 53506 45554 53518
rect 45502 53442 45554 53454
rect 46062 53506 46114 53518
rect 46062 53442 46114 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 1822 53170 1874 53182
rect 29038 53170 29090 53182
rect 23426 53118 23438 53170
rect 23490 53118 23502 53170
rect 1822 53106 1874 53118
rect 29038 53106 29090 53118
rect 29710 53170 29762 53182
rect 29710 53106 29762 53118
rect 3726 53058 3778 53070
rect 3726 52994 3778 53006
rect 3950 53058 4002 53070
rect 3950 52994 4002 53006
rect 6190 53058 6242 53070
rect 6190 52994 6242 53006
rect 14142 53058 14194 53070
rect 14142 52994 14194 53006
rect 18622 53058 18674 53070
rect 18622 52994 18674 53006
rect 28030 53058 28082 53070
rect 28030 52994 28082 53006
rect 28254 53058 28306 53070
rect 28254 52994 28306 53006
rect 30494 53058 30546 53070
rect 30494 52994 30546 53006
rect 31166 53058 31218 53070
rect 31166 52994 31218 53006
rect 42702 53058 42754 53070
rect 42702 52994 42754 53006
rect 43374 53058 43426 53070
rect 43374 52994 43426 53006
rect 9102 52946 9154 52958
rect 17054 52946 17106 52958
rect 31614 52946 31666 52958
rect 8530 52894 8542 52946
rect 8594 52894 8606 52946
rect 16482 52894 16494 52946
rect 16546 52894 16558 52946
rect 20514 52894 20526 52946
rect 20578 52894 20590 52946
rect 21074 52894 21086 52946
rect 21138 52894 21150 52946
rect 9102 52882 9154 52894
rect 17054 52882 17106 52894
rect 31614 52882 31666 52894
rect 3838 52834 3890 52846
rect 3838 52770 3890 52782
rect 4510 52834 4562 52846
rect 4510 52770 4562 52782
rect 9662 52834 9714 52846
rect 9662 52770 9714 52782
rect 10222 52834 10274 52846
rect 10222 52770 10274 52782
rect 10558 52834 10610 52846
rect 10558 52770 10610 52782
rect 12462 52834 12514 52846
rect 12462 52770 12514 52782
rect 17614 52834 17666 52846
rect 17614 52770 17666 52782
rect 18174 52834 18226 52846
rect 18174 52770 18226 52782
rect 19966 52834 20018 52846
rect 19966 52770 20018 52782
rect 24558 52834 24610 52846
rect 24558 52770 24610 52782
rect 27358 52834 27410 52846
rect 27358 52770 27410 52782
rect 29150 52834 29202 52846
rect 29150 52770 29202 52782
rect 29822 52834 29874 52846
rect 29822 52770 29874 52782
rect 39454 52834 39506 52846
rect 39454 52770 39506 52782
rect 40798 52834 40850 52846
rect 40798 52770 40850 52782
rect 41470 52834 41522 52846
rect 41470 52770 41522 52782
rect 43598 52834 43650 52846
rect 43598 52770 43650 52782
rect 44046 52834 44098 52846
rect 44046 52770 44098 52782
rect 5406 52722 5458 52734
rect 5406 52658 5458 52670
rect 13358 52722 13410 52734
rect 13358 52658 13410 52670
rect 24110 52722 24162 52734
rect 24110 52658 24162 52670
rect 27246 52722 27298 52734
rect 27246 52658 27298 52670
rect 27918 52722 27970 52734
rect 27918 52658 27970 52670
rect 30382 52722 30434 52734
rect 30382 52658 30434 52670
rect 31054 52722 31106 52734
rect 31054 52658 31106 52670
rect 43262 52722 43314 52734
rect 43262 52658 43314 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 31390 52386 31442 52398
rect 31390 52322 31442 52334
rect 51438 52386 51490 52398
rect 51438 52322 51490 52334
rect 11902 52274 11954 52286
rect 11902 52210 11954 52222
rect 20526 52274 20578 52286
rect 20526 52210 20578 52222
rect 21534 52274 21586 52286
rect 21534 52210 21586 52222
rect 28478 52274 28530 52286
rect 28478 52210 28530 52222
rect 29486 52274 29538 52286
rect 29486 52210 29538 52222
rect 30046 52274 30098 52286
rect 30046 52210 30098 52222
rect 30718 52274 30770 52286
rect 30718 52210 30770 52222
rect 31502 52274 31554 52286
rect 31502 52210 31554 52222
rect 52670 52274 52722 52286
rect 52670 52210 52722 52222
rect 7198 52162 7250 52174
rect 10894 52162 10946 52174
rect 10210 52110 10222 52162
rect 10274 52110 10286 52162
rect 7198 52098 7250 52110
rect 10894 52098 10946 52110
rect 11454 52162 11506 52174
rect 11454 52098 11506 52110
rect 16494 52162 16546 52174
rect 22094 52162 22146 52174
rect 16930 52110 16942 52162
rect 16994 52110 17006 52162
rect 16494 52098 16546 52110
rect 22094 52098 22146 52110
rect 27582 52162 27634 52174
rect 27582 52098 27634 52110
rect 28366 52162 28418 52174
rect 28366 52098 28418 52110
rect 51774 52162 51826 52174
rect 51774 52098 51826 52110
rect 52222 52162 52274 52174
rect 52222 52098 52274 52110
rect 53454 52162 53506 52174
rect 53454 52098 53506 52110
rect 53566 52162 53618 52174
rect 54114 52110 54126 52162
rect 54178 52110 54190 52162
rect 53566 52098 53618 52110
rect 19966 51938 20018 51950
rect 7970 51886 7982 51938
rect 8034 51886 8046 51938
rect 19170 51886 19182 51938
rect 19234 51886 19246 51938
rect 19966 51874 20018 51886
rect 31950 51938 32002 51950
rect 31950 51874 32002 51886
rect 51550 51938 51602 51950
rect 51550 51874 51602 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 40126 51602 40178 51614
rect 22642 51550 22654 51602
rect 22706 51550 22718 51602
rect 40126 51538 40178 51550
rect 53118 51602 53170 51614
rect 53118 51538 53170 51550
rect 3950 51490 4002 51502
rect 3950 51426 4002 51438
rect 4622 51490 4674 51502
rect 4622 51426 4674 51438
rect 18734 51490 18786 51502
rect 18734 51426 18786 51438
rect 11118 51378 11170 51390
rect 11118 51314 11170 51326
rect 19518 51378 19570 51390
rect 39902 51378 39954 51390
rect 40798 51378 40850 51390
rect 20178 51326 20190 51378
rect 20242 51326 20254 51378
rect 40226 51326 40238 51378
rect 40290 51326 40302 51378
rect 19518 51314 19570 51326
rect 39902 51314 39954 51326
rect 40798 51314 40850 51326
rect 43150 51378 43202 51390
rect 43474 51326 43486 51378
rect 43538 51326 43550 51378
rect 43150 51314 43202 51326
rect 5182 51266 5234 51278
rect 5182 51202 5234 51214
rect 11902 51266 11954 51278
rect 11902 51202 11954 51214
rect 18286 51266 18338 51278
rect 18286 51202 18338 51214
rect 23662 51266 23714 51278
rect 23662 51202 23714 51214
rect 38558 51266 38610 51278
rect 38558 51202 38610 51214
rect 39006 51266 39058 51278
rect 41582 51266 41634 51278
rect 40002 51214 40014 51266
rect 40066 51214 40078 51266
rect 39006 51202 39058 51214
rect 41582 51202 41634 51214
rect 42142 51266 42194 51278
rect 42142 51202 42194 51214
rect 42478 51266 42530 51278
rect 42478 51202 42530 51214
rect 43038 51266 43090 51278
rect 43038 51202 43090 51214
rect 3726 51154 3778 51166
rect 3726 51090 3778 51102
rect 4062 51154 4114 51166
rect 4062 51090 4114 51102
rect 4734 51154 4786 51166
rect 4734 51090 4786 51102
rect 23214 51154 23266 51166
rect 23214 51090 23266 51102
rect 40574 51154 40626 51166
rect 40574 51090 40626 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 40462 50818 40514 50830
rect 39106 50766 39118 50818
rect 39170 50815 39182 50818
rect 39778 50815 39790 50818
rect 39170 50769 39790 50815
rect 39170 50766 39182 50769
rect 39778 50766 39790 50769
rect 39842 50766 39854 50818
rect 40462 50754 40514 50766
rect 18622 50706 18674 50718
rect 18622 50642 18674 50654
rect 35534 50706 35586 50718
rect 40114 50654 40126 50706
rect 40178 50654 40190 50706
rect 35534 50642 35586 50654
rect 8206 50594 8258 50606
rect 19742 50594 19794 50606
rect 8642 50542 8654 50594
rect 8706 50542 8718 50594
rect 15026 50542 15038 50594
rect 15090 50542 15102 50594
rect 15586 50542 15598 50594
rect 15650 50542 15662 50594
rect 8206 50530 8258 50542
rect 19742 50530 19794 50542
rect 1822 50482 1874 50494
rect 1822 50418 1874 50430
rect 12238 50482 12290 50494
rect 12238 50418 12290 50430
rect 12686 50482 12738 50494
rect 12686 50418 12738 50430
rect 39454 50482 39506 50494
rect 39454 50418 39506 50430
rect 40238 50482 40290 50494
rect 40238 50418 40290 50430
rect 40910 50482 40962 50494
rect 40910 50418 40962 50430
rect 57262 50482 57314 50494
rect 57262 50418 57314 50430
rect 58046 50482 58098 50494
rect 58046 50418 58098 50430
rect 2158 50370 2210 50382
rect 11678 50370 11730 50382
rect 19182 50370 19234 50382
rect 11106 50318 11118 50370
rect 11170 50318 11182 50370
rect 18050 50318 18062 50370
rect 18114 50318 18126 50370
rect 2158 50306 2210 50318
rect 11678 50306 11730 50318
rect 19182 50306 19234 50318
rect 32398 50370 32450 50382
rect 32398 50306 32450 50318
rect 36094 50370 36146 50382
rect 36094 50306 36146 50318
rect 36654 50370 36706 50382
rect 36654 50306 36706 50318
rect 57710 50370 57762 50382
rect 57710 50306 57762 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 1822 50034 1874 50046
rect 43598 50034 43650 50046
rect 22082 49982 22094 50034
rect 22146 49982 22158 50034
rect 1822 49970 1874 49982
rect 43598 49970 43650 49982
rect 44270 50034 44322 50046
rect 44270 49970 44322 49982
rect 44942 50034 44994 50046
rect 44942 49970 44994 49982
rect 32174 49922 32226 49934
rect 12226 49870 12238 49922
rect 12290 49870 12302 49922
rect 32174 49858 32226 49870
rect 32622 49922 32674 49934
rect 32622 49858 32674 49870
rect 35870 49922 35922 49934
rect 35870 49858 35922 49870
rect 44494 49922 44546 49934
rect 44494 49858 44546 49870
rect 18958 49810 19010 49822
rect 36430 49810 36482 49822
rect 15026 49758 15038 49810
rect 15090 49758 15102 49810
rect 19618 49758 19630 49810
rect 19682 49758 19694 49810
rect 18958 49746 19010 49758
rect 36430 49746 36482 49758
rect 15598 49698 15650 49710
rect 15598 49634 15650 49646
rect 18510 49698 18562 49710
rect 18510 49634 18562 49646
rect 23102 49698 23154 49710
rect 23102 49634 23154 49646
rect 31502 49698 31554 49710
rect 31502 49634 31554 49646
rect 36878 49698 36930 49710
rect 36878 49634 36930 49646
rect 22654 49586 22706 49598
rect 22654 49522 22706 49534
rect 31390 49586 31442 49598
rect 31390 49522 31442 49534
rect 32062 49586 32114 49598
rect 32062 49522 32114 49534
rect 44158 49586 44210 49598
rect 44158 49522 44210 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 27682 49198 27694 49250
rect 27746 49247 27758 49250
rect 27906 49247 27918 49250
rect 27746 49201 27918 49247
rect 27746 49198 27758 49201
rect 27906 49198 27918 49201
rect 27970 49198 27982 49250
rect 11006 49138 11058 49150
rect 27918 49138 27970 49150
rect 18498 49086 18510 49138
rect 18562 49086 18574 49138
rect 11006 49074 11058 49086
rect 27918 49074 27970 49086
rect 31950 49138 32002 49150
rect 31950 49074 32002 49086
rect 32398 49138 32450 49150
rect 32398 49074 32450 49086
rect 35870 49138 35922 49150
rect 35870 49074 35922 49086
rect 10334 49026 10386 49038
rect 9762 48974 9774 49026
rect 9826 48974 9838 49026
rect 20514 48974 20526 49026
rect 20578 48974 20590 49026
rect 10334 48962 10386 48974
rect 31838 48914 31890 48926
rect 31838 48850 31890 48862
rect 6638 48802 6690 48814
rect 11342 48802 11394 48814
rect 7410 48750 7422 48802
rect 7474 48750 7486 48802
rect 6638 48738 6690 48750
rect 11342 48738 11394 48750
rect 21534 48802 21586 48814
rect 21534 48738 21586 48750
rect 36430 48802 36482 48814
rect 36430 48738 36482 48750
rect 37438 48802 37490 48814
rect 37438 48738 37490 48750
rect 47518 48802 47570 48814
rect 47518 48738 47570 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 4510 48466 4562 48478
rect 4510 48402 4562 48414
rect 10558 48466 10610 48478
rect 10558 48402 10610 48414
rect 12126 48466 12178 48478
rect 12126 48402 12178 48414
rect 46622 48466 46674 48478
rect 46622 48402 46674 48414
rect 47070 48466 47122 48478
rect 47070 48402 47122 48414
rect 3950 48354 4002 48366
rect 3950 48290 4002 48302
rect 27694 48354 27746 48366
rect 27694 48290 27746 48302
rect 48078 48354 48130 48366
rect 48078 48290 48130 48302
rect 48190 48354 48242 48366
rect 48190 48290 48242 48302
rect 37998 48242 38050 48254
rect 3042 48190 3054 48242
rect 3106 48190 3118 48242
rect 47842 48190 47854 48242
rect 47906 48190 47918 48242
rect 37998 48178 38050 48190
rect 28702 48130 28754 48142
rect 2034 48078 2046 48130
rect 2098 48078 2110 48130
rect 3938 48078 3950 48130
rect 4002 48078 4014 48130
rect 28702 48066 28754 48078
rect 29150 48130 29202 48142
rect 29150 48066 29202 48078
rect 38558 48130 38610 48142
rect 38558 48066 38610 48078
rect 3726 48018 3778 48030
rect 3726 47954 3778 47966
rect 27582 48018 27634 48030
rect 27582 47954 27634 47966
rect 28590 48018 28642 48030
rect 28590 47954 28642 47966
rect 37886 48018 37938 48030
rect 48626 47966 48638 48018
rect 48690 47966 48702 48018
rect 37886 47954 37938 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 19406 47570 19458 47582
rect 18386 47518 18398 47570
rect 18450 47518 18462 47570
rect 19406 47506 19458 47518
rect 26798 47570 26850 47582
rect 26798 47506 26850 47518
rect 27358 47570 27410 47582
rect 27358 47506 27410 47518
rect 46846 47570 46898 47582
rect 46846 47506 46898 47518
rect 47294 47570 47346 47582
rect 47294 47506 47346 47518
rect 49086 47570 49138 47582
rect 49086 47506 49138 47518
rect 8542 47458 8594 47470
rect 28030 47458 28082 47470
rect 8978 47406 8990 47458
rect 9042 47406 9054 47458
rect 14018 47406 14030 47458
rect 14082 47406 14094 47458
rect 8542 47394 8594 47406
rect 28030 47394 28082 47406
rect 48078 47458 48130 47470
rect 48078 47394 48130 47406
rect 48302 47458 48354 47470
rect 48302 47394 48354 47406
rect 48750 47458 48802 47470
rect 48750 47394 48802 47406
rect 28702 47346 28754 47358
rect 28702 47282 28754 47294
rect 3278 47234 3330 47246
rect 12014 47234 12066 47246
rect 11442 47182 11454 47234
rect 11506 47182 11518 47234
rect 3278 47170 3330 47182
rect 12014 47170 12066 47182
rect 12574 47234 12626 47246
rect 12574 47170 12626 47182
rect 27246 47234 27298 47246
rect 27246 47170 27298 47182
rect 27918 47234 27970 47246
rect 27918 47170 27970 47182
rect 28590 47234 28642 47246
rect 28590 47170 28642 47182
rect 29486 47234 29538 47246
rect 29486 47170 29538 47182
rect 48414 47234 48466 47246
rect 48414 47170 48466 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 4510 46898 4562 46910
rect 28254 46898 28306 46910
rect 23426 46846 23438 46898
rect 23490 46846 23502 46898
rect 4510 46834 4562 46846
rect 28254 46834 28306 46846
rect 28702 46898 28754 46910
rect 28702 46834 28754 46846
rect 29934 46898 29986 46910
rect 29934 46834 29986 46846
rect 43038 46898 43090 46910
rect 43038 46834 43090 46846
rect 4062 46786 4114 46798
rect 4062 46722 4114 46734
rect 27806 46786 27858 46798
rect 27806 46722 27858 46734
rect 29486 46786 29538 46798
rect 29486 46722 29538 46734
rect 20414 46674 20466 46686
rect 42926 46674 42978 46686
rect 3714 46622 3726 46674
rect 3778 46622 3790 46674
rect 21074 46622 21086 46674
rect 21138 46622 21150 46674
rect 20414 46610 20466 46622
rect 42926 46610 42978 46622
rect 43150 46674 43202 46686
rect 43150 46610 43202 46622
rect 43822 46674 43874 46686
rect 43822 46610 43874 46622
rect 47966 46674 48018 46686
rect 47966 46610 48018 46622
rect 3166 46562 3218 46574
rect 3166 46498 3218 46510
rect 9774 46562 9826 46574
rect 9774 46498 9826 46510
rect 12350 46562 12402 46574
rect 12350 46498 12402 46510
rect 19630 46562 19682 46574
rect 19630 46498 19682 46510
rect 20078 46562 20130 46574
rect 20078 46498 20130 46510
rect 24558 46562 24610 46574
rect 24558 46498 24610 46510
rect 29374 46562 29426 46574
rect 29374 46498 29426 46510
rect 32958 46562 33010 46574
rect 32958 46498 33010 46510
rect 33742 46562 33794 46574
rect 33742 46498 33794 46510
rect 34414 46562 34466 46574
rect 34414 46498 34466 46510
rect 34862 46562 34914 46574
rect 34862 46498 34914 46510
rect 37102 46562 37154 46574
rect 37102 46498 37154 46510
rect 37438 46562 37490 46574
rect 37438 46498 37490 46510
rect 41806 46562 41858 46574
rect 41806 46498 41858 46510
rect 42366 46562 42418 46574
rect 42366 46498 42418 46510
rect 43374 46562 43426 46574
rect 43374 46498 43426 46510
rect 47742 46562 47794 46574
rect 47742 46498 47794 46510
rect 48078 46562 48130 46574
rect 48078 46498 48130 46510
rect 48750 46562 48802 46574
rect 48750 46498 48802 46510
rect 3726 46450 3778 46462
rect 3726 46386 3778 46398
rect 24110 46450 24162 46462
rect 24110 46386 24162 46398
rect 27694 46450 27746 46462
rect 27694 46386 27746 46398
rect 33630 46450 33682 46462
rect 33630 46386 33682 46398
rect 34302 46450 34354 46462
rect 34302 46386 34354 46398
rect 43598 46450 43650 46462
rect 43598 46386 43650 46398
rect 47630 46450 47682 46462
rect 47630 46386 47682 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 35870 46114 35922 46126
rect 35870 46050 35922 46062
rect 38334 46114 38386 46126
rect 38334 46050 38386 46062
rect 11230 46002 11282 46014
rect 11230 45938 11282 45950
rect 31726 46002 31778 46014
rect 31726 45938 31778 45950
rect 32398 46002 32450 46014
rect 32398 45938 32450 45950
rect 35422 46002 35474 46014
rect 35422 45938 35474 45950
rect 10670 45890 10722 45902
rect 10098 45838 10110 45890
rect 10162 45838 10174 45890
rect 10670 45826 10722 45838
rect 11678 45890 11730 45902
rect 19630 45890 19682 45902
rect 19170 45838 19182 45890
rect 19234 45838 19246 45890
rect 11678 45826 11730 45838
rect 19630 45826 19682 45838
rect 30718 45890 30770 45902
rect 38558 45890 38610 45902
rect 35522 45838 35534 45890
rect 35586 45887 35598 45890
rect 35746 45887 35758 45890
rect 35586 45841 35758 45887
rect 35586 45838 35598 45841
rect 35746 45838 35758 45841
rect 35810 45838 35822 45890
rect 36194 45838 36206 45890
rect 36258 45838 36270 45890
rect 37986 45838 37998 45890
rect 38050 45838 38062 45890
rect 30718 45826 30770 45838
rect 38558 45826 38610 45838
rect 16158 45778 16210 45790
rect 16158 45714 16210 45726
rect 16942 45778 16994 45790
rect 16942 45714 16994 45726
rect 34078 45778 34130 45790
rect 34078 45714 34130 45726
rect 34526 45778 34578 45790
rect 34526 45714 34578 45726
rect 6974 45666 7026 45678
rect 20414 45666 20466 45678
rect 7746 45614 7758 45666
rect 7810 45614 7822 45666
rect 6974 45602 7026 45614
rect 20414 45602 20466 45614
rect 20862 45666 20914 45678
rect 20862 45602 20914 45614
rect 28702 45666 28754 45678
rect 28702 45602 28754 45614
rect 30606 45666 30658 45678
rect 30606 45602 30658 45614
rect 31166 45666 31218 45678
rect 31166 45602 31218 45614
rect 33966 45666 34018 45678
rect 33966 45602 34018 45614
rect 35982 45666 36034 45678
rect 35982 45602 36034 45614
rect 36654 45666 36706 45678
rect 36654 45602 36706 45614
rect 37662 45666 37714 45678
rect 37662 45602 37714 45614
rect 37774 45666 37826 45678
rect 37774 45602 37826 45614
rect 37886 45666 37938 45678
rect 37886 45602 37938 45614
rect 39006 45666 39058 45678
rect 39006 45602 39058 45614
rect 40350 45666 40402 45678
rect 40350 45602 40402 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2158 45330 2210 45342
rect 27582 45330 27634 45342
rect 23314 45278 23326 45330
rect 23378 45278 23390 45330
rect 2158 45266 2210 45278
rect 27582 45266 27634 45278
rect 29934 45330 29986 45342
rect 29934 45266 29986 45278
rect 30718 45330 30770 45342
rect 30718 45266 30770 45278
rect 32622 45330 32674 45342
rect 32622 45266 32674 45278
rect 39902 45330 39954 45342
rect 39902 45266 39954 45278
rect 40798 45330 40850 45342
rect 40798 45266 40850 45278
rect 6190 45218 6242 45230
rect 6190 45154 6242 45166
rect 31502 45218 31554 45230
rect 31502 45154 31554 45166
rect 32174 45218 32226 45230
rect 32174 45154 32226 45166
rect 37326 45218 37378 45230
rect 37326 45154 37378 45166
rect 38222 45218 38274 45230
rect 38222 45154 38274 45166
rect 39790 45218 39842 45230
rect 39790 45154 39842 45166
rect 40686 45218 40738 45230
rect 40686 45154 40738 45166
rect 1822 45106 1874 45118
rect 8878 45106 8930 45118
rect 8530 45054 8542 45106
rect 8594 45054 8606 45106
rect 1822 45042 1874 45054
rect 8878 45042 8930 45054
rect 11230 45106 11282 45118
rect 11230 45042 11282 45054
rect 20190 45106 20242 45118
rect 29262 45106 29314 45118
rect 20738 45054 20750 45106
rect 20802 45054 20814 45106
rect 20190 45042 20242 45054
rect 29262 45042 29314 45054
rect 29710 45106 29762 45118
rect 29710 45042 29762 45054
rect 30158 45106 30210 45118
rect 36978 45054 36990 45106
rect 37042 45054 37054 45106
rect 30158 45042 30210 45054
rect 9774 44994 9826 45006
rect 9774 44930 9826 44942
rect 10110 44994 10162 45006
rect 10110 44930 10162 44942
rect 10782 44994 10834 45006
rect 10782 44930 10834 44942
rect 19742 44994 19794 45006
rect 19742 44930 19794 44942
rect 24334 44994 24386 45006
rect 24334 44930 24386 44942
rect 27918 44994 27970 45006
rect 27918 44930 27970 44942
rect 28590 44994 28642 45006
rect 37214 44994 37266 45006
rect 30034 44942 30046 44994
rect 30098 44942 30110 44994
rect 28590 44930 28642 44942
rect 37214 44930 37266 44942
rect 37774 44994 37826 45006
rect 37774 44930 37826 44942
rect 40014 44994 40066 45006
rect 40014 44930 40066 44942
rect 41582 44994 41634 45006
rect 41582 44930 41634 44942
rect 5406 44882 5458 44894
rect 5406 44818 5458 44830
rect 23886 44882 23938 44894
rect 23886 44818 23938 44830
rect 28478 44882 28530 44894
rect 28478 44818 28530 44830
rect 29486 44882 29538 44894
rect 29486 44818 29538 44830
rect 31390 44882 31442 44894
rect 31390 44818 31442 44830
rect 32062 44882 32114 44894
rect 32062 44818 32114 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 30158 44546 30210 44558
rect 40002 44494 40014 44546
rect 40066 44543 40078 44546
rect 40226 44543 40238 44546
rect 40066 44497 40238 44543
rect 40066 44494 40078 44497
rect 40226 44494 40238 44497
rect 40290 44494 40302 44546
rect 30158 44482 30210 44494
rect 1822 44434 1874 44446
rect 1822 44370 1874 44382
rect 28814 44434 28866 44446
rect 28814 44370 28866 44382
rect 30270 44434 30322 44446
rect 30270 44370 30322 44382
rect 31166 44434 31218 44446
rect 31166 44370 31218 44382
rect 31950 44434 32002 44446
rect 31950 44370 32002 44382
rect 33518 44434 33570 44446
rect 33518 44370 33570 44382
rect 11118 44322 11170 44334
rect 10546 44270 10558 44322
rect 10610 44270 10622 44322
rect 11118 44258 11170 44270
rect 12126 44322 12178 44334
rect 12126 44258 12178 44270
rect 15038 44322 15090 44334
rect 31054 44322 31106 44334
rect 15362 44270 15374 44322
rect 15426 44270 15438 44322
rect 15038 44258 15090 44270
rect 31054 44258 31106 44270
rect 19294 44210 19346 44222
rect 19294 44146 19346 44158
rect 32510 44210 32562 44222
rect 32510 44146 32562 44158
rect 58046 44210 58098 44222
rect 58046 44146 58098 44158
rect 7422 44098 7474 44110
rect 11678 44098 11730 44110
rect 8194 44046 8206 44098
rect 8258 44046 8270 44098
rect 7422 44034 7474 44046
rect 11678 44034 11730 44046
rect 14366 44098 14418 44110
rect 18510 44098 18562 44110
rect 17938 44046 17950 44098
rect 18002 44046 18014 44098
rect 14366 44034 14418 44046
rect 18510 44034 18562 44046
rect 18846 44098 18898 44110
rect 18846 44034 18898 44046
rect 31838 44098 31890 44110
rect 31838 44034 31890 44046
rect 32622 44098 32674 44110
rect 32622 44034 32674 44046
rect 33070 44098 33122 44110
rect 33070 44034 33122 44046
rect 40238 44098 40290 44110
rect 40238 44034 40290 44046
rect 57262 44098 57314 44110
rect 57262 44034 57314 44046
rect 57710 44098 57762 44110
rect 57710 44034 57762 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 30606 43762 30658 43774
rect 6178 43710 6190 43762
rect 6242 43710 6254 43762
rect 16146 43710 16158 43762
rect 16210 43710 16222 43762
rect 23426 43710 23438 43762
rect 23490 43710 23502 43762
rect 30606 43698 30658 43710
rect 32510 43762 32562 43774
rect 32510 43698 32562 43710
rect 36766 43762 36818 43774
rect 36766 43698 36818 43710
rect 10222 43650 10274 43662
rect 10222 43586 10274 43598
rect 17726 43650 17778 43662
rect 17726 43586 17778 43598
rect 24334 43650 24386 43662
rect 24334 43586 24386 43598
rect 24894 43650 24946 43662
rect 24894 43586 24946 43598
rect 31614 43650 31666 43662
rect 31614 43586 31666 43598
rect 32062 43650 32114 43662
rect 32062 43586 32114 43598
rect 33966 43650 34018 43662
rect 33966 43586 34018 43598
rect 36878 43650 36930 43662
rect 36878 43586 36930 43598
rect 8878 43538 8930 43550
rect 8530 43486 8542 43538
rect 8594 43486 8606 43538
rect 8878 43474 8930 43486
rect 13022 43538 13074 43550
rect 20302 43538 20354 43550
rect 36654 43538 36706 43550
rect 13570 43486 13582 43538
rect 13634 43486 13646 43538
rect 20962 43486 20974 43538
rect 21026 43486 21038 43538
rect 35074 43486 35086 43538
rect 35138 43486 35150 43538
rect 13022 43474 13074 43486
rect 20302 43474 20354 43486
rect 36654 43474 36706 43486
rect 9662 43426 9714 43438
rect 9662 43362 9714 43374
rect 10782 43426 10834 43438
rect 10782 43362 10834 43374
rect 11342 43426 11394 43438
rect 11342 43362 11394 43374
rect 12126 43426 12178 43438
rect 12126 43362 12178 43374
rect 12686 43426 12738 43438
rect 12686 43362 12738 43374
rect 19854 43426 19906 43438
rect 19854 43362 19906 43374
rect 33854 43426 33906 43438
rect 33854 43362 33906 43374
rect 35534 43426 35586 43438
rect 35534 43362 35586 43374
rect 35982 43426 36034 43438
rect 35982 43362 36034 43374
rect 37102 43426 37154 43438
rect 37102 43362 37154 43374
rect 5406 43314 5458 43326
rect 5406 43250 5458 43262
rect 16718 43314 16770 43326
rect 16718 43250 16770 43262
rect 23998 43314 24050 43326
rect 23998 43250 24050 43262
rect 31502 43314 31554 43326
rect 31502 43250 31554 43262
rect 34750 43314 34802 43326
rect 34750 43250 34802 43262
rect 35086 43314 35138 43326
rect 35086 43250 35138 43262
rect 37326 43314 37378 43326
rect 37326 43250 37378 43262
rect 37550 43314 37602 43326
rect 37550 43250 37602 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 10670 42866 10722 42878
rect 10670 42802 10722 42814
rect 12910 42866 12962 42878
rect 12910 42802 12962 42814
rect 34638 42866 34690 42878
rect 34638 42802 34690 42814
rect 6638 42754 6690 42766
rect 13582 42754 13634 42766
rect 17614 42754 17666 42766
rect 7074 42702 7086 42754
rect 7138 42702 7150 42754
rect 14242 42702 14254 42754
rect 14306 42702 14318 42754
rect 6638 42690 6690 42702
rect 13582 42690 13634 42702
rect 17614 42690 17666 42702
rect 33742 42754 33794 42766
rect 34178 42702 34190 42754
rect 34242 42702 34254 42754
rect 33742 42690 33794 42702
rect 16494 42642 16546 42654
rect 16494 42578 16546 42590
rect 18062 42642 18114 42654
rect 18062 42578 18114 42590
rect 45614 42642 45666 42654
rect 45614 42578 45666 42590
rect 10110 42530 10162 42542
rect 9538 42478 9550 42530
rect 9602 42478 9614 42530
rect 10110 42466 10162 42478
rect 11118 42530 11170 42542
rect 11118 42466 11170 42478
rect 17278 42530 17330 42542
rect 17278 42466 17330 42478
rect 36206 42530 36258 42542
rect 36206 42466 36258 42478
rect 45502 42530 45554 42542
rect 45502 42466 45554 42478
rect 46062 42530 46114 42542
rect 46062 42466 46114 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 2158 42194 2210 42206
rect 23202 42142 23214 42194
rect 23266 42142 23278 42194
rect 2158 42130 2210 42142
rect 10658 42030 10670 42082
rect 10722 42030 10734 42082
rect 1822 41970 1874 41982
rect 20078 41970 20130 41982
rect 24670 41970 24722 41982
rect 15026 41918 15038 41970
rect 15090 41918 15102 41970
rect 20738 41918 20750 41970
rect 20802 41918 20814 41970
rect 1822 41906 1874 41918
rect 20078 41906 20130 41918
rect 24670 41906 24722 41918
rect 15486 41858 15538 41870
rect 15486 41794 15538 41806
rect 19630 41858 19682 41870
rect 19630 41794 19682 41806
rect 24222 41858 24274 41870
rect 24222 41794 24274 41806
rect 23774 41746 23826 41758
rect 23774 41682 23826 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 1822 41298 1874 41310
rect 1822 41234 1874 41246
rect 11006 41298 11058 41310
rect 11006 41234 11058 41246
rect 28814 41298 28866 41310
rect 28814 41234 28866 41246
rect 34190 41298 34242 41310
rect 34190 41234 34242 41246
rect 35534 41298 35586 41310
rect 35534 41234 35586 41246
rect 36430 41298 36482 41310
rect 36430 41234 36482 41246
rect 37886 41298 37938 41310
rect 37886 41234 37938 41246
rect 42814 41298 42866 41310
rect 42814 41234 42866 41246
rect 10334 41186 10386 41198
rect 21534 41186 21586 41198
rect 9762 41134 9774 41186
rect 9826 41134 9838 41186
rect 16706 41134 16718 41186
rect 16770 41134 16782 41186
rect 10334 41122 10386 41134
rect 21534 41122 21586 41134
rect 42142 41186 42194 41198
rect 42142 41122 42194 41134
rect 42590 41186 42642 41198
rect 42590 41122 42642 41134
rect 42926 41186 42978 41198
rect 42926 41122 42978 41134
rect 29598 41074 29650 41086
rect 17378 41022 17390 41074
rect 17442 41022 17454 41074
rect 29598 41010 29650 41022
rect 29822 41074 29874 41086
rect 29822 41010 29874 41022
rect 33630 41074 33682 41086
rect 33630 41010 33682 41022
rect 33742 41074 33794 41086
rect 33742 41010 33794 41022
rect 35982 41074 36034 41086
rect 35982 41010 36034 41022
rect 41806 41074 41858 41086
rect 41806 41010 41858 41022
rect 41918 41074 41970 41086
rect 41918 41010 41970 41022
rect 43262 41074 43314 41086
rect 43262 41010 43314 41022
rect 57262 41074 57314 41086
rect 57262 41010 57314 41022
rect 58046 41074 58098 41086
rect 58046 41010 58098 41022
rect 6638 40962 6690 40974
rect 11342 40962 11394 40974
rect 7410 40910 7422 40962
rect 7474 40910 7486 40962
rect 6638 40898 6690 40910
rect 11342 40898 11394 40910
rect 29710 40962 29762 40974
rect 29710 40898 29762 40910
rect 33406 40962 33458 40974
rect 33406 40898 33458 40910
rect 35086 40962 35138 40974
rect 35086 40898 35138 40910
rect 37550 40962 37602 40974
rect 37550 40898 37602 40910
rect 43822 40962 43874 40974
rect 43822 40898 43874 40910
rect 57710 40962 57762 40974
rect 57710 40898 57762 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 22766 40626 22818 40638
rect 22194 40574 22206 40626
rect 22258 40574 22270 40626
rect 22766 40562 22818 40574
rect 23662 40626 23714 40638
rect 23662 40562 23714 40574
rect 25902 40626 25954 40638
rect 25902 40562 25954 40574
rect 26350 40626 26402 40638
rect 26350 40562 26402 40574
rect 26798 40626 26850 40638
rect 26798 40562 26850 40574
rect 28366 40626 28418 40638
rect 28366 40562 28418 40574
rect 30046 40626 30098 40638
rect 30046 40562 30098 40574
rect 31390 40626 31442 40638
rect 31390 40562 31442 40574
rect 32062 40626 32114 40638
rect 32062 40562 32114 40574
rect 32622 40626 32674 40638
rect 32622 40562 32674 40574
rect 34862 40626 34914 40638
rect 34862 40562 34914 40574
rect 35758 40626 35810 40638
rect 35758 40562 35810 40574
rect 35870 40626 35922 40638
rect 35870 40562 35922 40574
rect 40686 40626 40738 40638
rect 40686 40562 40738 40574
rect 42478 40626 42530 40638
rect 42478 40562 42530 40574
rect 42702 40626 42754 40638
rect 42702 40562 42754 40574
rect 10558 40514 10610 40526
rect 10558 40450 10610 40462
rect 18622 40514 18674 40526
rect 31054 40514 31106 40526
rect 27458 40462 27470 40514
rect 27522 40462 27534 40514
rect 27794 40462 27806 40514
rect 27858 40462 27870 40514
rect 18622 40450 18674 40462
rect 31054 40450 31106 40462
rect 31166 40514 31218 40526
rect 40014 40514 40066 40526
rect 38770 40462 38782 40514
rect 38834 40462 38846 40514
rect 31166 40450 31218 40462
rect 40014 40450 40066 40462
rect 47630 40514 47682 40526
rect 47630 40450 47682 40462
rect 19070 40402 19122 40414
rect 23214 40402 23266 40414
rect 30494 40402 30546 40414
rect 19730 40350 19742 40402
rect 19794 40350 19806 40402
rect 27906 40350 27918 40402
rect 27970 40350 27982 40402
rect 19070 40338 19122 40350
rect 23214 40338 23266 40350
rect 30494 40338 30546 40350
rect 34302 40402 34354 40414
rect 34302 40338 34354 40350
rect 35982 40402 36034 40414
rect 35982 40338 36034 40350
rect 36206 40402 36258 40414
rect 41470 40402 41522 40414
rect 37538 40350 37550 40402
rect 37602 40350 37614 40402
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 38546 40350 38558 40402
rect 38610 40350 38622 40402
rect 36206 40338 36258 40350
rect 41470 40338 41522 40350
rect 42142 40402 42194 40414
rect 42142 40338 42194 40350
rect 43150 40402 43202 40414
rect 43150 40338 43202 40350
rect 47518 40402 47570 40414
rect 47518 40338 47570 40350
rect 47854 40402 47906 40414
rect 47854 40338 47906 40350
rect 27358 40290 27410 40302
rect 27358 40226 27410 40238
rect 31838 40290 31890 40302
rect 35086 40290 35138 40302
rect 32050 40238 32062 40290
rect 32114 40238 32126 40290
rect 31838 40226 31890 40238
rect 35086 40226 35138 40238
rect 36654 40290 36706 40302
rect 40238 40290 40290 40302
rect 39890 40238 39902 40290
rect 39954 40238 39966 40290
rect 36654 40226 36706 40238
rect 40238 40226 40290 40238
rect 48190 40290 48242 40302
rect 48190 40226 48242 40238
rect 34750 40178 34802 40190
rect 34750 40114 34802 40126
rect 36430 40178 36482 40190
rect 36430 40114 36482 40126
rect 37214 40178 37266 40190
rect 37214 40114 37266 40126
rect 42814 40178 42866 40190
rect 42814 40114 42866 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 20078 39842 20130 39854
rect 20078 39778 20130 39790
rect 33854 39842 33906 39854
rect 33854 39778 33906 39790
rect 40574 39842 40626 39854
rect 40574 39778 40626 39790
rect 20638 39730 20690 39742
rect 20638 39666 20690 39678
rect 27246 39730 27298 39742
rect 27246 39666 27298 39678
rect 28702 39730 28754 39742
rect 28702 39666 28754 39678
rect 37438 39730 37490 39742
rect 37438 39666 37490 39678
rect 38334 39730 38386 39742
rect 38334 39666 38386 39678
rect 41134 39730 41186 39742
rect 41134 39666 41186 39678
rect 42030 39730 42082 39742
rect 42030 39666 42082 39678
rect 42478 39730 42530 39742
rect 42478 39666 42530 39678
rect 16606 39618 16658 39630
rect 21534 39618 21586 39630
rect 17042 39566 17054 39618
rect 17106 39566 17118 39618
rect 16606 39554 16658 39566
rect 21534 39554 21586 39566
rect 28366 39618 28418 39630
rect 28366 39554 28418 39566
rect 28478 39618 28530 39630
rect 28478 39554 28530 39566
rect 31838 39618 31890 39630
rect 31838 39554 31890 39566
rect 35086 39618 35138 39630
rect 35086 39554 35138 39566
rect 35646 39618 35698 39630
rect 35646 39554 35698 39566
rect 38110 39618 38162 39630
rect 38110 39554 38162 39566
rect 38558 39618 38610 39630
rect 38558 39554 38610 39566
rect 39902 39618 39954 39630
rect 39902 39554 39954 39566
rect 40462 39618 40514 39630
rect 40462 39554 40514 39566
rect 47518 39618 47570 39630
rect 47518 39554 47570 39566
rect 48302 39618 48354 39630
rect 48302 39554 48354 39566
rect 28814 39506 28866 39518
rect 28814 39442 28866 39454
rect 31278 39506 31330 39518
rect 31278 39442 31330 39454
rect 31502 39506 31554 39518
rect 31502 39442 31554 39454
rect 32286 39506 32338 39518
rect 32286 39442 32338 39454
rect 33742 39506 33794 39518
rect 33742 39442 33794 39454
rect 34750 39506 34802 39518
rect 34750 39442 34802 39454
rect 34862 39506 34914 39518
rect 34862 39442 34914 39454
rect 36206 39506 36258 39518
rect 36206 39442 36258 39454
rect 38782 39506 38834 39518
rect 38782 39442 38834 39454
rect 39230 39506 39282 39518
rect 39230 39442 39282 39454
rect 40574 39506 40626 39518
rect 40574 39442 40626 39454
rect 47294 39506 47346 39518
rect 47294 39442 47346 39454
rect 48750 39506 48802 39518
rect 48750 39442 48802 39454
rect 48974 39506 49026 39518
rect 48974 39442 49026 39454
rect 26350 39394 26402 39406
rect 19506 39342 19518 39394
rect 19570 39342 19582 39394
rect 26350 39330 26402 39342
rect 26798 39394 26850 39406
rect 26798 39330 26850 39342
rect 27806 39394 27858 39406
rect 27806 39330 27858 39342
rect 31614 39394 31666 39406
rect 31614 39330 31666 39342
rect 33182 39394 33234 39406
rect 33182 39330 33234 39342
rect 35758 39394 35810 39406
rect 35758 39330 35810 39342
rect 35982 39394 36034 39406
rect 35982 39330 36034 39342
rect 36318 39394 36370 39406
rect 36318 39330 36370 39342
rect 36654 39394 36706 39406
rect 36654 39330 36706 39342
rect 41582 39394 41634 39406
rect 41582 39330 41634 39342
rect 46734 39394 46786 39406
rect 48526 39394 48578 39406
rect 47842 39342 47854 39394
rect 47906 39342 47918 39394
rect 46734 39330 46786 39342
rect 48526 39330 48578 39342
rect 49422 39394 49474 39406
rect 49422 39330 49474 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 2158 39058 2210 39070
rect 2158 38994 2210 39006
rect 20414 39058 20466 39070
rect 20414 38994 20466 39006
rect 27582 39058 27634 39070
rect 27582 38994 27634 39006
rect 30942 39058 30994 39070
rect 30942 38994 30994 39006
rect 34974 39058 35026 39070
rect 34974 38994 35026 39006
rect 35422 39058 35474 39070
rect 35422 38994 35474 39006
rect 35758 39058 35810 39070
rect 35758 38994 35810 39006
rect 36430 39058 36482 39070
rect 44158 39058 44210 39070
rect 39218 39006 39230 39058
rect 39282 39006 39294 39058
rect 36430 38994 36482 39006
rect 44158 38994 44210 39006
rect 45278 39058 45330 39070
rect 45278 38994 45330 39006
rect 45502 39058 45554 39070
rect 45502 38994 45554 39006
rect 46622 39058 46674 39070
rect 46622 38994 46674 39006
rect 27022 38946 27074 38958
rect 50766 38946 50818 38958
rect 39106 38894 39118 38946
rect 39170 38894 39182 38946
rect 40562 38894 40574 38946
rect 40626 38894 40638 38946
rect 27022 38882 27074 38894
rect 50766 38882 50818 38894
rect 51326 38946 51378 38958
rect 51326 38882 51378 38894
rect 1822 38834 1874 38846
rect 1822 38770 1874 38782
rect 38558 38834 38610 38846
rect 45390 38834 45442 38846
rect 38994 38782 39006 38834
rect 39058 38782 39070 38834
rect 40674 38782 40686 38834
rect 40738 38782 40750 38834
rect 38558 38770 38610 38782
rect 45390 38770 45442 38782
rect 45950 38834 46002 38846
rect 45950 38770 46002 38782
rect 3838 38722 3890 38734
rect 3838 38658 3890 38670
rect 4398 38722 4450 38734
rect 4398 38658 4450 38670
rect 13134 38722 13186 38734
rect 13134 38658 13186 38670
rect 13694 38722 13746 38734
rect 13694 38658 13746 38670
rect 14702 38722 14754 38734
rect 14702 38658 14754 38670
rect 15150 38722 15202 38734
rect 15150 38658 15202 38670
rect 34414 38722 34466 38734
rect 34414 38658 34466 38670
rect 41582 38722 41634 38734
rect 41582 38658 41634 38670
rect 41918 38722 41970 38734
rect 41918 38658 41970 38670
rect 44606 38722 44658 38734
rect 44606 38658 44658 38670
rect 45726 38722 45778 38734
rect 45726 38658 45778 38670
rect 3950 38610 4002 38622
rect 3950 38546 4002 38558
rect 26910 38610 26962 38622
rect 26910 38546 26962 38558
rect 46174 38610 46226 38622
rect 46174 38546 46226 38558
rect 50878 38610 50930 38622
rect 50878 38546 50930 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 26574 38274 26626 38286
rect 26574 38210 26626 38222
rect 1822 38162 1874 38174
rect 1822 38098 1874 38110
rect 12014 38162 12066 38174
rect 12014 38098 12066 38110
rect 24558 38162 24610 38174
rect 24558 38098 24610 38110
rect 34414 38162 34466 38174
rect 41694 38162 41746 38174
rect 35074 38110 35086 38162
rect 35138 38110 35150 38162
rect 41122 38110 41134 38162
rect 41186 38110 41198 38162
rect 34414 38098 34466 38110
rect 41694 38098 41746 38110
rect 14590 38050 14642 38062
rect 14242 37998 14254 38050
rect 14306 37998 14318 38050
rect 14590 37986 14642 37998
rect 25566 38050 25618 38062
rect 30830 38050 30882 38062
rect 26114 37998 26126 38050
rect 26178 37998 26190 38050
rect 25566 37986 25618 37998
rect 30830 37986 30882 37998
rect 31166 38050 31218 38062
rect 31166 37986 31218 37998
rect 31502 38050 31554 38062
rect 31502 37986 31554 37998
rect 32846 38050 32898 38062
rect 32846 37986 32898 37998
rect 33518 38050 33570 38062
rect 33518 37986 33570 37998
rect 33966 38050 34018 38062
rect 39454 38050 39506 38062
rect 35298 37998 35310 38050
rect 35362 37998 35374 38050
rect 33966 37986 34018 37998
rect 39454 37986 39506 37998
rect 39790 38050 39842 38062
rect 42142 38050 42194 38062
rect 40898 37998 40910 38050
rect 40962 37998 40974 38050
rect 39790 37986 39842 37998
rect 42142 37986 42194 37998
rect 12910 37938 12962 37950
rect 12910 37874 12962 37886
rect 14030 37938 14082 37950
rect 14030 37874 14082 37886
rect 15150 37938 15202 37950
rect 25902 37938 25954 37950
rect 25666 37886 25678 37938
rect 25730 37886 25742 37938
rect 15150 37874 15202 37886
rect 25902 37874 25954 37886
rect 30158 37938 30210 37950
rect 30158 37874 30210 37886
rect 30382 37938 30434 37950
rect 30382 37874 30434 37886
rect 35982 37938 36034 37950
rect 35982 37874 36034 37886
rect 36654 37938 36706 37950
rect 36654 37874 36706 37886
rect 39118 37938 39170 37950
rect 39118 37874 39170 37886
rect 40238 37938 40290 37950
rect 40238 37874 40290 37886
rect 58046 37938 58098 37950
rect 58046 37874 58098 37886
rect 12686 37826 12738 37838
rect 12686 37762 12738 37774
rect 12798 37826 12850 37838
rect 12798 37762 12850 37774
rect 13918 37826 13970 37838
rect 13918 37762 13970 37774
rect 15038 37826 15090 37838
rect 15038 37762 15090 37774
rect 15598 37826 15650 37838
rect 15598 37762 15650 37774
rect 18510 37826 18562 37838
rect 18510 37762 18562 37774
rect 19070 37826 19122 37838
rect 19070 37762 19122 37774
rect 24110 37826 24162 37838
rect 24110 37762 24162 37774
rect 25006 37826 25058 37838
rect 25006 37762 25058 37774
rect 26910 37826 26962 37838
rect 26910 37762 26962 37774
rect 27358 37826 27410 37838
rect 27358 37762 27410 37774
rect 30606 37826 30658 37838
rect 30606 37762 30658 37774
rect 31390 37826 31442 37838
rect 31390 37762 31442 37774
rect 31950 37826 32002 37838
rect 31950 37762 32002 37774
rect 32398 37826 32450 37838
rect 32398 37762 32450 37774
rect 32958 37826 33010 37838
rect 32958 37762 33010 37774
rect 33182 37826 33234 37838
rect 33182 37762 33234 37774
rect 36542 37826 36594 37838
rect 36542 37762 36594 37774
rect 39454 37826 39506 37838
rect 39454 37762 39506 37774
rect 57262 37826 57314 37838
rect 57262 37762 57314 37774
rect 57710 37826 57762 37838
rect 57710 37762 57762 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 10894 37490 10946 37502
rect 10894 37426 10946 37438
rect 13358 37490 13410 37502
rect 13358 37426 13410 37438
rect 16942 37490 16994 37502
rect 16942 37426 16994 37438
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 20526 37490 20578 37502
rect 32622 37490 32674 37502
rect 27346 37438 27358 37490
rect 27410 37438 27422 37490
rect 20526 37426 20578 37438
rect 32622 37426 32674 37438
rect 36206 37490 36258 37502
rect 36206 37426 36258 37438
rect 12014 37378 12066 37390
rect 12014 37314 12066 37326
rect 17726 37378 17778 37390
rect 17726 37314 17778 37326
rect 25006 37378 25058 37390
rect 25006 37314 25058 37326
rect 25790 37378 25842 37390
rect 31502 37378 31554 37390
rect 27234 37326 27246 37378
rect 27298 37326 27310 37378
rect 30930 37326 30942 37378
rect 30994 37326 31006 37378
rect 25790 37314 25842 37326
rect 31502 37314 31554 37326
rect 40462 37378 40514 37390
rect 40462 37314 40514 37326
rect 40686 37378 40738 37390
rect 40686 37314 40738 37326
rect 12574 37266 12626 37278
rect 12574 37202 12626 37214
rect 12798 37266 12850 37278
rect 12798 37202 12850 37214
rect 13246 37266 13298 37278
rect 13246 37202 13298 37214
rect 13470 37266 13522 37278
rect 13470 37202 13522 37214
rect 19294 37266 19346 37278
rect 19294 37202 19346 37214
rect 19742 37266 19794 37278
rect 19742 37202 19794 37214
rect 19966 37266 20018 37278
rect 19966 37202 20018 37214
rect 20974 37266 21026 37278
rect 20974 37202 21026 37214
rect 25678 37266 25730 37278
rect 25678 37202 25730 37214
rect 28814 37266 28866 37278
rect 41470 37266 41522 37278
rect 29138 37214 29150 37266
rect 29202 37214 29214 37266
rect 28814 37202 28866 37214
rect 41470 37202 41522 37214
rect 49646 37266 49698 37278
rect 49970 37214 49982 37266
rect 50034 37214 50046 37266
rect 49646 37202 49698 37214
rect 5070 37154 5122 37166
rect 5070 37090 5122 37102
rect 8766 37154 8818 37166
rect 8766 37090 8818 37102
rect 11454 37154 11506 37166
rect 11454 37090 11506 37102
rect 13022 37154 13074 37166
rect 13022 37090 13074 37102
rect 14030 37154 14082 37166
rect 14030 37090 14082 37102
rect 14478 37154 14530 37166
rect 14478 37090 14530 37102
rect 14926 37154 14978 37166
rect 14926 37090 14978 37102
rect 15374 37154 15426 37166
rect 15374 37090 15426 37102
rect 16494 37154 16546 37166
rect 16494 37090 16546 37102
rect 18510 37154 18562 37166
rect 18510 37090 18562 37102
rect 19518 37154 19570 37166
rect 19518 37090 19570 37102
rect 26574 37154 26626 37166
rect 26574 37090 26626 37102
rect 39790 37154 39842 37166
rect 39790 37090 39842 37102
rect 40574 37154 40626 37166
rect 40574 37090 40626 37102
rect 49534 37154 49586 37166
rect 49534 37090 49586 37102
rect 50990 37154 51042 37166
rect 50990 37090 51042 37102
rect 11902 37042 11954 37054
rect 11902 36978 11954 36990
rect 17838 37042 17890 37054
rect 17838 36978 17890 36990
rect 19070 37042 19122 37054
rect 19070 36978 19122 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 3838 36706 3890 36718
rect 3838 36642 3890 36654
rect 31054 36706 31106 36718
rect 31054 36642 31106 36654
rect 34078 36706 34130 36718
rect 34078 36642 34130 36654
rect 41358 36706 41410 36718
rect 41358 36642 41410 36654
rect 42478 36706 42530 36718
rect 42478 36642 42530 36654
rect 49534 36706 49586 36718
rect 49534 36642 49586 36654
rect 4062 36594 4114 36606
rect 5630 36594 5682 36606
rect 11454 36594 11506 36606
rect 13694 36594 13746 36606
rect 16942 36594 16994 36606
rect 4498 36542 4510 36594
rect 4562 36542 4574 36594
rect 8082 36542 8094 36594
rect 8146 36542 8158 36594
rect 8866 36542 8878 36594
rect 8930 36542 8942 36594
rect 12674 36542 12686 36594
rect 12738 36542 12750 36594
rect 14578 36542 14590 36594
rect 14642 36542 14654 36594
rect 4062 36530 4114 36542
rect 5630 36530 5682 36542
rect 11454 36530 11506 36542
rect 13694 36530 13746 36542
rect 16942 36530 16994 36542
rect 17390 36594 17442 36606
rect 19854 36594 19906 36606
rect 19058 36542 19070 36594
rect 19122 36542 19134 36594
rect 17390 36530 17442 36542
rect 19854 36530 19906 36542
rect 20414 36594 20466 36606
rect 27134 36594 27186 36606
rect 32286 36594 32338 36606
rect 24882 36542 24894 36594
rect 24946 36542 24958 36594
rect 30482 36542 30494 36594
rect 30546 36542 30558 36594
rect 20414 36530 20466 36542
rect 27134 36530 27186 36542
rect 32286 36530 32338 36542
rect 32734 36594 32786 36606
rect 32734 36530 32786 36542
rect 34414 36594 34466 36606
rect 34414 36530 34466 36542
rect 34862 36594 34914 36606
rect 41582 36594 41634 36606
rect 42926 36594 42978 36606
rect 40786 36542 40798 36594
rect 40850 36542 40862 36594
rect 42130 36542 42142 36594
rect 42194 36542 42206 36594
rect 34862 36530 34914 36542
rect 41582 36530 41634 36542
rect 42926 36530 42978 36542
rect 43486 36594 43538 36606
rect 43486 36530 43538 36542
rect 6414 36482 6466 36494
rect 4386 36430 4398 36482
rect 4450 36430 4462 36482
rect 6414 36418 6466 36430
rect 7310 36482 7362 36494
rect 7310 36418 7362 36430
rect 7534 36482 7586 36494
rect 8206 36482 8258 36494
rect 7858 36430 7870 36482
rect 7922 36430 7934 36482
rect 7534 36418 7586 36430
rect 8206 36418 8258 36430
rect 11902 36482 11954 36494
rect 11902 36418 11954 36430
rect 12126 36482 12178 36494
rect 19182 36482 19234 36494
rect 12450 36430 12462 36482
rect 12514 36430 12526 36482
rect 14130 36430 14142 36482
rect 14194 36430 14206 36482
rect 12126 36418 12178 36430
rect 19182 36418 19234 36430
rect 19406 36482 19458 36494
rect 19406 36418 19458 36430
rect 19630 36482 19682 36494
rect 19630 36418 19682 36430
rect 25230 36482 25282 36494
rect 25230 36418 25282 36430
rect 25454 36482 25506 36494
rect 25454 36418 25506 36430
rect 25678 36482 25730 36494
rect 25678 36418 25730 36430
rect 30606 36482 30658 36494
rect 31278 36482 31330 36494
rect 30706 36430 30718 36482
rect 30770 36430 30782 36482
rect 30606 36418 30658 36430
rect 31278 36418 31330 36430
rect 32174 36482 32226 36494
rect 32174 36418 32226 36430
rect 33518 36482 33570 36494
rect 41134 36482 41186 36494
rect 34066 36430 34078 36482
rect 34130 36430 34142 36482
rect 33518 36418 33570 36430
rect 41134 36418 41186 36430
rect 1822 36370 1874 36382
rect 1822 36306 1874 36318
rect 8990 36370 9042 36382
rect 8990 36306 9042 36318
rect 9214 36370 9266 36382
rect 9214 36306 9266 36318
rect 12798 36370 12850 36382
rect 12798 36306 12850 36318
rect 15934 36370 15986 36382
rect 15934 36306 15986 36318
rect 16158 36370 16210 36382
rect 16158 36306 16210 36318
rect 18286 36370 18338 36382
rect 18286 36306 18338 36318
rect 23550 36370 23602 36382
rect 23550 36306 23602 36318
rect 24110 36370 24162 36382
rect 24110 36306 24162 36318
rect 40014 36370 40066 36382
rect 40014 36306 40066 36318
rect 42254 36370 42306 36382
rect 42254 36306 42306 36318
rect 2158 36258 2210 36270
rect 2158 36194 2210 36206
rect 4510 36258 4562 36270
rect 4510 36194 4562 36206
rect 4734 36258 4786 36270
rect 4734 36194 4786 36206
rect 6862 36258 6914 36270
rect 6862 36194 6914 36206
rect 7982 36258 8034 36270
rect 7982 36194 8034 36206
rect 9774 36258 9826 36270
rect 9774 36194 9826 36206
rect 10110 36258 10162 36270
rect 10110 36194 10162 36206
rect 10558 36258 10610 36270
rect 10558 36194 10610 36206
rect 12574 36258 12626 36270
rect 12574 36194 12626 36206
rect 15374 36258 15426 36270
rect 15374 36194 15426 36206
rect 16046 36258 16098 36270
rect 16046 36194 16098 36206
rect 16830 36258 16882 36270
rect 16830 36194 16882 36206
rect 17838 36258 17890 36270
rect 17838 36194 17890 36206
rect 18958 36258 19010 36270
rect 18958 36194 19010 36206
rect 22878 36258 22930 36270
rect 22878 36194 22930 36206
rect 23438 36258 23490 36270
rect 23438 36194 23490 36206
rect 24782 36258 24834 36270
rect 24782 36194 24834 36206
rect 25006 36258 25058 36270
rect 25006 36194 25058 36206
rect 26238 36258 26290 36270
rect 26238 36194 26290 36206
rect 26574 36258 26626 36270
rect 26574 36194 26626 36206
rect 29710 36258 29762 36270
rect 29710 36194 29762 36206
rect 30382 36258 30434 36270
rect 30382 36194 30434 36206
rect 39566 36258 39618 36270
rect 39566 36194 39618 36206
rect 40686 36258 40738 36270
rect 40686 36194 40738 36206
rect 40910 36258 40962 36270
rect 40910 36194 40962 36206
rect 49310 36258 49362 36270
rect 49310 36194 49362 36206
rect 49422 36258 49474 36270
rect 49422 36194 49474 36206
rect 49982 36258 50034 36270
rect 49982 36194 50034 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 5294 35922 5346 35934
rect 5294 35858 5346 35870
rect 8206 35922 8258 35934
rect 8206 35858 8258 35870
rect 14142 35922 14194 35934
rect 14142 35858 14194 35870
rect 14702 35922 14754 35934
rect 14702 35858 14754 35870
rect 16158 35922 16210 35934
rect 17838 35922 17890 35934
rect 17154 35870 17166 35922
rect 17218 35870 17230 35922
rect 16158 35858 16210 35870
rect 1710 35810 1762 35822
rect 1710 35746 1762 35758
rect 8766 35810 8818 35822
rect 8766 35746 8818 35758
rect 8878 35810 8930 35822
rect 12910 35810 12962 35822
rect 9762 35758 9774 35810
rect 9826 35758 9838 35810
rect 8878 35746 8930 35758
rect 12910 35746 12962 35758
rect 14254 35810 14306 35822
rect 14254 35746 14306 35758
rect 15374 35810 15426 35822
rect 15374 35746 15426 35758
rect 9102 35698 9154 35710
rect 16046 35698 16098 35710
rect 10098 35646 10110 35698
rect 10162 35646 10174 35698
rect 9102 35634 9154 35646
rect 16046 35634 16098 35646
rect 16270 35698 16322 35710
rect 16270 35634 16322 35646
rect 16494 35698 16546 35710
rect 16494 35634 16546 35646
rect 16718 35698 16770 35710
rect 16718 35634 16770 35646
rect 16942 35698 16994 35710
rect 16942 35634 16994 35646
rect 11342 35586 11394 35598
rect 10434 35534 10446 35586
rect 10498 35534 10510 35586
rect 11342 35522 11394 35534
rect 11790 35586 11842 35598
rect 11790 35522 11842 35534
rect 13358 35586 13410 35598
rect 13358 35522 13410 35534
rect 17169 35474 17215 35870
rect 17838 35858 17890 35870
rect 18734 35922 18786 35934
rect 18734 35858 18786 35870
rect 20078 35922 20130 35934
rect 20078 35858 20130 35870
rect 32846 35922 32898 35934
rect 32846 35858 32898 35870
rect 35982 35922 36034 35934
rect 35982 35858 36034 35870
rect 39678 35922 39730 35934
rect 39678 35858 39730 35870
rect 44718 35922 44770 35934
rect 44718 35858 44770 35870
rect 45166 35922 45218 35934
rect 45166 35858 45218 35870
rect 45950 35922 46002 35934
rect 45950 35858 46002 35870
rect 46062 35922 46114 35934
rect 46062 35858 46114 35870
rect 18286 35810 18338 35822
rect 18286 35746 18338 35758
rect 29710 35810 29762 35822
rect 35646 35810 35698 35822
rect 33618 35758 33630 35810
rect 33682 35758 33694 35810
rect 35074 35758 35086 35810
rect 35138 35758 35150 35810
rect 29710 35746 29762 35758
rect 35646 35746 35698 35758
rect 35758 35810 35810 35822
rect 35758 35746 35810 35758
rect 38222 35810 38274 35822
rect 38222 35746 38274 35758
rect 39566 35810 39618 35822
rect 39566 35746 39618 35758
rect 45838 35810 45890 35822
rect 45838 35746 45890 35758
rect 47294 35810 47346 35822
rect 47294 35746 47346 35758
rect 49534 35810 49586 35822
rect 49534 35746 49586 35758
rect 19294 35698 19346 35710
rect 19966 35698 20018 35710
rect 19842 35646 19854 35698
rect 19906 35646 19918 35698
rect 19294 35634 19346 35646
rect 19966 35634 20018 35646
rect 20190 35698 20242 35710
rect 20190 35634 20242 35646
rect 32398 35698 32450 35710
rect 39790 35698 39842 35710
rect 33730 35646 33742 35698
rect 33794 35646 33806 35698
rect 34402 35646 34414 35698
rect 34466 35646 34478 35698
rect 34962 35646 34974 35698
rect 35026 35646 35038 35698
rect 32398 35634 32450 35646
rect 39790 35634 39842 35646
rect 46286 35698 46338 35710
rect 46286 35634 46338 35646
rect 46510 35698 46562 35710
rect 46510 35634 46562 35646
rect 50094 35698 50146 35710
rect 50094 35634 50146 35646
rect 50878 35698 50930 35710
rect 50878 35634 50930 35646
rect 51886 35698 51938 35710
rect 51886 35634 51938 35646
rect 31502 35586 31554 35598
rect 31502 35522 31554 35534
rect 36318 35586 36370 35598
rect 36318 35522 36370 35534
rect 38670 35586 38722 35598
rect 38670 35522 38722 35534
rect 40014 35586 40066 35598
rect 40014 35522 40066 35534
rect 41806 35586 41858 35598
rect 51314 35534 51326 35586
rect 51378 35534 51390 35586
rect 41806 35522 41858 35534
rect 19518 35474 19570 35486
rect 17154 35422 17166 35474
rect 17218 35422 17230 35474
rect 19518 35410 19570 35422
rect 40238 35474 40290 35486
rect 40238 35410 40290 35422
rect 40462 35474 40514 35486
rect 40462 35410 40514 35422
rect 46734 35474 46786 35486
rect 46734 35410 46786 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 19406 35138 19458 35150
rect 24782 35138 24834 35150
rect 23650 35086 23662 35138
rect 23714 35135 23726 35138
rect 24546 35135 24558 35138
rect 23714 35089 24558 35135
rect 23714 35086 23726 35089
rect 24546 35086 24558 35089
rect 24610 35086 24622 35138
rect 19406 35074 19458 35086
rect 24782 35074 24834 35086
rect 29598 35138 29650 35150
rect 29598 35074 29650 35086
rect 8990 35026 9042 35038
rect 8990 34962 9042 34974
rect 12238 35026 12290 35038
rect 15934 35026 15986 35038
rect 15138 34974 15150 35026
rect 15202 34974 15214 35026
rect 12238 34962 12290 34974
rect 15934 34962 15986 34974
rect 16942 35026 16994 35038
rect 16942 34962 16994 34974
rect 21870 35026 21922 35038
rect 21870 34962 21922 34974
rect 22430 35026 22482 35038
rect 22430 34962 22482 34974
rect 22990 35026 23042 35038
rect 26686 35026 26738 35038
rect 25442 34974 25454 35026
rect 25506 34974 25518 35026
rect 22990 34962 23042 34974
rect 26686 34962 26738 34974
rect 33294 35026 33346 35038
rect 33294 34962 33346 34974
rect 35646 35026 35698 35038
rect 35646 34962 35698 34974
rect 44718 35026 44770 35038
rect 44718 34962 44770 34974
rect 46062 35026 46114 35038
rect 46062 34962 46114 34974
rect 56254 35026 56306 35038
rect 57810 34974 57822 35026
rect 57874 34974 57886 35026
rect 56254 34962 56306 34974
rect 11678 34914 11730 34926
rect 17614 34914 17666 34926
rect 25006 34914 25058 34926
rect 15474 34862 15486 34914
rect 15538 34862 15550 34914
rect 17938 34862 17950 34914
rect 18002 34862 18014 34914
rect 22082 34862 22094 34914
rect 22146 34862 22158 34914
rect 11678 34850 11730 34862
rect 17614 34850 17666 34862
rect 25006 34850 25058 34862
rect 25230 34914 25282 34926
rect 25230 34850 25282 34862
rect 26350 34914 26402 34926
rect 26350 34850 26402 34862
rect 34526 34914 34578 34926
rect 34526 34850 34578 34862
rect 34862 34914 34914 34926
rect 34862 34850 34914 34862
rect 35086 34914 35138 34926
rect 35086 34850 35138 34862
rect 40238 34914 40290 34926
rect 40238 34850 40290 34862
rect 40462 34914 40514 34926
rect 45826 34862 45838 34914
rect 45890 34862 45902 34914
rect 56802 34862 56814 34914
rect 56866 34862 56878 34914
rect 40462 34850 40514 34862
rect 9550 34802 9602 34814
rect 9550 34738 9602 34750
rect 10222 34802 10274 34814
rect 10222 34738 10274 34750
rect 10558 34802 10610 34814
rect 10558 34738 10610 34750
rect 10782 34802 10834 34814
rect 10782 34738 10834 34750
rect 18510 34802 18562 34814
rect 18510 34738 18562 34750
rect 19070 34802 19122 34814
rect 19070 34738 19122 34750
rect 25454 34802 25506 34814
rect 25454 34738 25506 34750
rect 29710 34802 29762 34814
rect 29710 34738 29762 34750
rect 46174 34802 46226 34814
rect 46174 34738 46226 34750
rect 9662 34690 9714 34702
rect 9662 34626 9714 34638
rect 10334 34690 10386 34702
rect 10334 34626 10386 34638
rect 19294 34690 19346 34702
rect 19294 34626 19346 34638
rect 19854 34690 19906 34702
rect 19854 34626 19906 34638
rect 20414 34690 20466 34702
rect 20414 34626 20466 34638
rect 20862 34690 20914 34702
rect 20862 34626 20914 34638
rect 21758 34690 21810 34702
rect 21758 34626 21810 34638
rect 21982 34690 22034 34702
rect 21982 34626 22034 34638
rect 23326 34690 23378 34702
rect 23326 34626 23378 34638
rect 23774 34690 23826 34702
rect 23774 34626 23826 34638
rect 24222 34690 24274 34702
rect 24222 34626 24274 34638
rect 25678 34690 25730 34702
rect 25678 34626 25730 34638
rect 30158 34690 30210 34702
rect 30158 34626 30210 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 36094 34690 36146 34702
rect 36094 34626 36146 34638
rect 39118 34690 39170 34702
rect 46622 34690 46674 34702
rect 39890 34638 39902 34690
rect 39954 34638 39966 34690
rect 39118 34626 39170 34638
rect 46622 34626 46674 34638
rect 50318 34690 50370 34702
rect 50318 34626 50370 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 8542 34354 8594 34366
rect 8542 34290 8594 34302
rect 10558 34354 10610 34366
rect 10558 34290 10610 34302
rect 34414 34354 34466 34366
rect 34414 34290 34466 34302
rect 34526 34354 34578 34366
rect 34526 34290 34578 34302
rect 36094 34354 36146 34366
rect 36094 34290 36146 34302
rect 36542 34354 36594 34366
rect 36542 34290 36594 34302
rect 37438 34354 37490 34366
rect 37438 34290 37490 34302
rect 45166 34354 45218 34366
rect 45166 34290 45218 34302
rect 45838 34354 45890 34366
rect 45838 34290 45890 34302
rect 45950 34354 46002 34366
rect 45950 34290 46002 34302
rect 4734 34242 4786 34254
rect 4734 34178 4786 34190
rect 7982 34242 8034 34254
rect 7982 34178 8034 34190
rect 8094 34242 8146 34254
rect 8094 34178 8146 34190
rect 10446 34242 10498 34254
rect 36754 34190 36766 34242
rect 36818 34190 36830 34242
rect 10446 34178 10498 34190
rect 9998 34130 10050 34142
rect 5058 34078 5070 34130
rect 5122 34078 5134 34130
rect 9998 34066 10050 34078
rect 10670 34130 10722 34142
rect 10670 34066 10722 34078
rect 11230 34130 11282 34142
rect 11230 34066 11282 34078
rect 34638 34130 34690 34142
rect 34638 34066 34690 34078
rect 35086 34130 35138 34142
rect 35086 34066 35138 34078
rect 5518 34018 5570 34030
rect 4946 33966 4958 34018
rect 5010 33966 5022 34018
rect 5518 33954 5570 33966
rect 9774 34018 9826 34030
rect 9774 33954 9826 33966
rect 10222 34018 10274 34030
rect 10222 33954 10274 33966
rect 11678 34018 11730 34030
rect 11678 33954 11730 33966
rect 19854 34018 19906 34030
rect 19854 33954 19906 33966
rect 20414 34018 20466 34030
rect 20414 33954 20466 33966
rect 26574 34018 26626 34030
rect 26574 33954 26626 33966
rect 27022 34018 27074 34030
rect 27022 33954 27074 33966
rect 33854 34018 33906 34030
rect 33854 33954 33906 33966
rect 35646 34018 35698 34030
rect 35646 33954 35698 33966
rect 19966 33906 20018 33918
rect 36194 33854 36206 33906
rect 36258 33903 36270 33906
rect 36769 33903 36815 34190
rect 36990 34018 37042 34030
rect 36990 33954 37042 33966
rect 37886 34018 37938 34030
rect 37886 33954 37938 33966
rect 46622 34018 46674 34030
rect 46622 33954 46674 33966
rect 46062 33906 46114 33918
rect 36258 33857 36815 33903
rect 36258 33854 36270 33857
rect 37426 33854 37438 33906
rect 37490 33903 37502 33906
rect 37986 33903 37998 33906
rect 37490 33857 37998 33903
rect 37490 33854 37502 33857
rect 37986 33854 37998 33857
rect 38050 33854 38062 33906
rect 46274 33854 46286 33906
rect 46338 33903 46350 33906
rect 46610 33903 46622 33906
rect 46338 33857 46622 33903
rect 46338 33854 46350 33857
rect 46610 33854 46622 33857
rect 46674 33854 46686 33906
rect 19966 33842 20018 33854
rect 46062 33842 46114 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 26462 33570 26514 33582
rect 26462 33506 26514 33518
rect 32622 33570 32674 33582
rect 32622 33506 32674 33518
rect 34750 33570 34802 33582
rect 34750 33506 34802 33518
rect 34974 33570 35026 33582
rect 34974 33506 35026 33518
rect 35198 33570 35250 33582
rect 35198 33506 35250 33518
rect 38334 33570 38386 33582
rect 38334 33506 38386 33518
rect 11454 33458 11506 33470
rect 11454 33394 11506 33406
rect 11902 33458 11954 33470
rect 11902 33394 11954 33406
rect 17278 33458 17330 33470
rect 17278 33394 17330 33406
rect 23998 33458 24050 33470
rect 23998 33394 24050 33406
rect 24446 33458 24498 33470
rect 24446 33394 24498 33406
rect 25454 33458 25506 33470
rect 25454 33394 25506 33406
rect 30270 33458 30322 33470
rect 30270 33394 30322 33406
rect 36318 33458 36370 33470
rect 42030 33458 42082 33470
rect 40002 33406 40014 33458
rect 40066 33406 40078 33458
rect 36318 33394 36370 33406
rect 42030 33394 42082 33406
rect 42478 33458 42530 33470
rect 42478 33394 42530 33406
rect 49534 33458 49586 33470
rect 49534 33394 49586 33406
rect 16158 33346 16210 33358
rect 16158 33282 16210 33294
rect 16718 33346 16770 33358
rect 16718 33282 16770 33294
rect 25790 33346 25842 33358
rect 35422 33346 35474 33358
rect 26114 33294 26126 33346
rect 26178 33294 26190 33346
rect 25790 33282 25842 33294
rect 35422 33282 35474 33294
rect 36094 33346 36146 33358
rect 36094 33282 36146 33294
rect 36766 33346 36818 33358
rect 38558 33346 38610 33358
rect 37986 33294 37998 33346
rect 38050 33294 38062 33346
rect 36766 33282 36818 33294
rect 38558 33282 38610 33294
rect 41918 33346 41970 33358
rect 41918 33282 41970 33294
rect 26798 33234 26850 33246
rect 25554 33182 25566 33234
rect 25618 33182 25630 33234
rect 26798 33170 26850 33182
rect 27022 33234 27074 33246
rect 27022 33170 27074 33182
rect 27134 33234 27186 33246
rect 27134 33170 27186 33182
rect 27806 33234 27858 33246
rect 27806 33170 27858 33182
rect 28254 33234 28306 33246
rect 28254 33170 28306 33182
rect 29598 33234 29650 33246
rect 29598 33170 29650 33182
rect 29710 33234 29762 33246
rect 29710 33170 29762 33182
rect 32286 33234 32338 33246
rect 32286 33170 32338 33182
rect 36542 33234 36594 33246
rect 36542 33170 36594 33182
rect 25006 33122 25058 33134
rect 25006 33058 25058 33070
rect 27694 33122 27746 33134
rect 27694 33058 27746 33070
rect 28926 33122 28978 33134
rect 28926 33058 28978 33070
rect 29934 33122 29986 33134
rect 29934 33058 29986 33070
rect 31726 33122 31778 33134
rect 31726 33058 31778 33070
rect 32510 33122 32562 33134
rect 32510 33058 32562 33070
rect 33070 33122 33122 33134
rect 33070 33058 33122 33070
rect 34302 33122 34354 33134
rect 34302 33058 34354 33070
rect 37662 33122 37714 33134
rect 37662 33058 37714 33070
rect 37774 33122 37826 33134
rect 37774 33058 37826 33070
rect 37886 33122 37938 33134
rect 37886 33058 37938 33070
rect 39006 33122 39058 33134
rect 39006 33058 39058 33070
rect 39566 33122 39618 33134
rect 39566 33058 39618 33070
rect 50094 33122 50146 33134
rect 50094 33058 50146 33070
rect 50542 33122 50594 33134
rect 50542 33058 50594 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 3502 32786 3554 32798
rect 3502 32722 3554 32734
rect 9998 32786 10050 32798
rect 9998 32722 10050 32734
rect 11454 32786 11506 32798
rect 11454 32722 11506 32734
rect 12238 32786 12290 32798
rect 12238 32722 12290 32734
rect 21646 32786 21698 32798
rect 21646 32722 21698 32734
rect 22542 32786 22594 32798
rect 22542 32722 22594 32734
rect 26350 32786 26402 32798
rect 26350 32722 26402 32734
rect 27246 32786 27298 32798
rect 27246 32722 27298 32734
rect 27358 32786 27410 32798
rect 27358 32722 27410 32734
rect 27470 32786 27522 32798
rect 27470 32722 27522 32734
rect 28590 32786 28642 32798
rect 28590 32722 28642 32734
rect 33966 32786 34018 32798
rect 33966 32722 34018 32734
rect 34526 32786 34578 32798
rect 34526 32722 34578 32734
rect 34750 32786 34802 32798
rect 34750 32722 34802 32734
rect 35534 32786 35586 32798
rect 35534 32722 35586 32734
rect 37214 32786 37266 32798
rect 37214 32722 37266 32734
rect 38222 32786 38274 32798
rect 38222 32722 38274 32734
rect 38894 32786 38946 32798
rect 38894 32722 38946 32734
rect 39566 32786 39618 32798
rect 39566 32722 39618 32734
rect 11566 32674 11618 32686
rect 11566 32610 11618 32622
rect 12462 32674 12514 32686
rect 12462 32610 12514 32622
rect 35310 32674 35362 32686
rect 35310 32610 35362 32622
rect 37326 32674 37378 32686
rect 37326 32610 37378 32622
rect 42702 32674 42754 32686
rect 42702 32610 42754 32622
rect 9886 32562 9938 32574
rect 3042 32510 3054 32562
rect 3106 32510 3118 32562
rect 9886 32498 9938 32510
rect 10110 32562 10162 32574
rect 10110 32498 10162 32510
rect 10334 32562 10386 32574
rect 10334 32498 10386 32510
rect 10782 32562 10834 32574
rect 10782 32498 10834 32510
rect 11230 32562 11282 32574
rect 11230 32498 11282 32510
rect 12014 32562 12066 32574
rect 12014 32498 12066 32510
rect 12574 32562 12626 32574
rect 12574 32498 12626 32510
rect 21422 32562 21474 32574
rect 21422 32498 21474 32510
rect 21758 32562 21810 32574
rect 21758 32498 21810 32510
rect 22206 32562 22258 32574
rect 22206 32498 22258 32510
rect 22654 32562 22706 32574
rect 22654 32498 22706 32510
rect 22878 32562 22930 32574
rect 22878 32498 22930 32510
rect 26014 32562 26066 32574
rect 26014 32498 26066 32510
rect 26238 32562 26290 32574
rect 26238 32498 26290 32510
rect 26686 32562 26738 32574
rect 34414 32562 34466 32574
rect 27570 32510 27582 32562
rect 27634 32510 27646 32562
rect 26686 32498 26738 32510
rect 34414 32498 34466 32510
rect 35198 32562 35250 32574
rect 35198 32498 35250 32510
rect 42142 32562 42194 32574
rect 42142 32498 42194 32510
rect 13134 32450 13186 32462
rect 2034 32398 2046 32450
rect 2098 32398 2110 32450
rect 13134 32386 13186 32398
rect 23326 32450 23378 32462
rect 23326 32386 23378 32398
rect 23774 32450 23826 32462
rect 23774 32386 23826 32398
rect 24894 32450 24946 32462
rect 24894 32386 24946 32398
rect 35870 32450 35922 32462
rect 35870 32386 35922 32398
rect 36318 32450 36370 32462
rect 40126 32450 40178 32462
rect 38098 32398 38110 32450
rect 38162 32398 38174 32450
rect 36318 32386 36370 32398
rect 40126 32386 40178 32398
rect 40686 32450 40738 32462
rect 40686 32386 40738 32398
rect 10558 32338 10610 32350
rect 10558 32274 10610 32286
rect 27918 32338 27970 32350
rect 27918 32274 27970 32286
rect 28142 32338 28194 32350
rect 28142 32274 28194 32286
rect 38446 32338 38498 32350
rect 38446 32274 38498 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 11006 31890 11058 31902
rect 11006 31826 11058 31838
rect 16046 31890 16098 31902
rect 16046 31826 16098 31838
rect 17166 31890 17218 31902
rect 17166 31826 17218 31838
rect 17502 31890 17554 31902
rect 26910 31890 26962 31902
rect 23650 31838 23662 31890
rect 23714 31838 23726 31890
rect 17502 31826 17554 31838
rect 26910 31826 26962 31838
rect 27246 31890 27298 31902
rect 35758 31890 35810 31902
rect 39902 31890 39954 31902
rect 30482 31838 30494 31890
rect 30546 31838 30558 31890
rect 39218 31838 39230 31890
rect 39282 31838 39294 31890
rect 27246 31826 27298 31838
rect 35758 31826 35810 31838
rect 39902 31826 39954 31838
rect 36878 31778 36930 31790
rect 36878 31714 36930 31726
rect 38110 31778 38162 31790
rect 41806 31778 41858 31790
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 39106 31726 39118 31778
rect 39170 31726 39182 31778
rect 38110 31714 38162 31726
rect 41806 31714 41858 31726
rect 11902 31666 11954 31678
rect 11902 31602 11954 31614
rect 16606 31666 16658 31678
rect 16606 31602 16658 31614
rect 17054 31666 17106 31678
rect 17054 31602 17106 31614
rect 23886 31666 23938 31678
rect 23886 31602 23938 31614
rect 30830 31666 30882 31678
rect 30830 31602 30882 31614
rect 37886 31666 37938 31678
rect 37886 31602 37938 31614
rect 37998 31666 38050 31678
rect 37998 31602 38050 31614
rect 39454 31666 39506 31678
rect 39454 31602 39506 31614
rect 41246 31666 41298 31678
rect 41246 31602 41298 31614
rect 11678 31554 11730 31566
rect 11678 31490 11730 31502
rect 11790 31554 11842 31566
rect 11790 31490 11842 31502
rect 12350 31554 12402 31566
rect 12350 31490 12402 31502
rect 16830 31554 16882 31566
rect 16830 31490 16882 31502
rect 18062 31554 18114 31566
rect 18062 31490 18114 31502
rect 21982 31554 22034 31566
rect 21982 31490 22034 31502
rect 23662 31554 23714 31566
rect 23662 31490 23714 31502
rect 24334 31554 24386 31566
rect 24334 31490 24386 31502
rect 24782 31554 24834 31566
rect 24782 31490 24834 31502
rect 30606 31554 30658 31566
rect 30606 31490 30658 31502
rect 31278 31554 31330 31566
rect 31278 31490 31330 31502
rect 31726 31554 31778 31566
rect 31726 31490 31778 31502
rect 34078 31554 34130 31566
rect 34078 31490 34130 31502
rect 40350 31554 40402 31566
rect 40350 31490 40402 31502
rect 41358 31554 41410 31566
rect 41358 31490 41410 31502
rect 58046 31554 58098 31566
rect 58046 31490 58098 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 10446 31218 10498 31230
rect 10446 31154 10498 31166
rect 10894 31218 10946 31230
rect 10894 31154 10946 31166
rect 29486 31218 29538 31230
rect 29486 31154 29538 31166
rect 39902 31218 39954 31230
rect 39902 31154 39954 31166
rect 40014 31218 40066 31230
rect 40014 31154 40066 31166
rect 40574 31218 40626 31230
rect 40574 31154 40626 31166
rect 12014 31106 12066 31118
rect 12014 31042 12066 31054
rect 12126 31106 12178 31118
rect 12126 31042 12178 31054
rect 12686 31106 12738 31118
rect 12686 31042 12738 31054
rect 11342 30994 11394 31006
rect 5506 30942 5518 30994
rect 5570 30942 5582 30994
rect 13122 30942 13134 30994
rect 13186 30942 13198 30994
rect 28914 30942 28926 30994
rect 28978 30942 28990 30994
rect 11342 30930 11394 30942
rect 4734 30882 4786 30894
rect 4734 30818 4786 30830
rect 5182 30882 5234 30894
rect 5182 30818 5234 30830
rect 5966 30882 6018 30894
rect 19070 30882 19122 30894
rect 13010 30830 13022 30882
rect 13074 30830 13086 30882
rect 5966 30818 6018 30830
rect 19070 30818 19122 30830
rect 28142 30882 28194 30894
rect 28142 30818 28194 30830
rect 28702 30882 28754 30894
rect 28702 30818 28754 30830
rect 37438 30882 37490 30894
rect 37438 30818 37490 30830
rect 40126 30882 40178 30894
rect 40126 30818 40178 30830
rect 41582 30882 41634 30894
rect 41582 30818 41634 30830
rect 5518 30770 5570 30782
rect 5518 30706 5570 30718
rect 12014 30770 12066 30782
rect 12014 30706 12066 30718
rect 28590 30770 28642 30782
rect 28590 30706 28642 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 8654 30434 8706 30446
rect 8654 30370 8706 30382
rect 9214 30434 9266 30446
rect 9214 30370 9266 30382
rect 9438 30434 9490 30446
rect 9438 30370 9490 30382
rect 19182 30434 19234 30446
rect 19182 30370 19234 30382
rect 32062 30434 32114 30446
rect 32062 30370 32114 30382
rect 5742 30322 5794 30334
rect 17726 30322 17778 30334
rect 6066 30270 6078 30322
rect 6130 30270 6142 30322
rect 5742 30258 5794 30270
rect 17726 30258 17778 30270
rect 6526 30210 6578 30222
rect 6526 30146 6578 30158
rect 9662 30210 9714 30222
rect 9662 30146 9714 30158
rect 9886 30210 9938 30222
rect 9886 30146 9938 30158
rect 9998 30210 10050 30222
rect 9998 30146 10050 30158
rect 10670 30210 10722 30222
rect 10670 30146 10722 30158
rect 12350 30210 12402 30222
rect 12350 30146 12402 30158
rect 12798 30210 12850 30222
rect 12798 30146 12850 30158
rect 13582 30210 13634 30222
rect 13582 30146 13634 30158
rect 13918 30210 13970 30222
rect 13918 30146 13970 30158
rect 14366 30210 14418 30222
rect 14366 30146 14418 30158
rect 16046 30210 16098 30222
rect 16046 30146 16098 30158
rect 17166 30210 17218 30222
rect 17166 30146 17218 30158
rect 17950 30210 18002 30222
rect 18622 30210 18674 30222
rect 19854 30210 19906 30222
rect 18274 30158 18286 30210
rect 18338 30158 18350 30210
rect 19618 30158 19630 30210
rect 19682 30158 19694 30210
rect 17950 30146 18002 30158
rect 18622 30146 18674 30158
rect 19854 30146 19906 30158
rect 20190 30210 20242 30222
rect 20190 30146 20242 30158
rect 21646 30210 21698 30222
rect 21646 30146 21698 30158
rect 1822 30098 1874 30110
rect 1822 30034 1874 30046
rect 2158 30098 2210 30110
rect 2158 30034 2210 30046
rect 5966 30098 6018 30110
rect 5966 30034 6018 30046
rect 8318 30098 8370 30110
rect 8318 30034 8370 30046
rect 8542 30098 8594 30110
rect 8542 30034 8594 30046
rect 10110 30098 10162 30110
rect 10110 30034 10162 30046
rect 12238 30098 12290 30110
rect 12238 30034 12290 30046
rect 13806 30098 13858 30110
rect 13806 30034 13858 30046
rect 14926 30098 14978 30110
rect 14926 30034 14978 30046
rect 15486 30098 15538 30110
rect 15486 30034 15538 30046
rect 19966 30098 20018 30110
rect 19966 30034 20018 30046
rect 20862 30098 20914 30110
rect 20862 30034 20914 30046
rect 32622 30098 32674 30110
rect 32622 30034 32674 30046
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 11342 29986 11394 29998
rect 11342 29922 11394 29934
rect 16830 29986 16882 29998
rect 16830 29922 16882 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 18510 29986 18562 29998
rect 18510 29922 18562 29934
rect 31166 29986 31218 29998
rect 31166 29922 31218 29934
rect 31614 29986 31666 29998
rect 31614 29922 31666 29934
rect 32174 29986 32226 29998
rect 32174 29922 32226 29934
rect 32398 29986 32450 29998
rect 32398 29922 32450 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 1822 29650 1874 29662
rect 1822 29586 1874 29598
rect 8990 29650 9042 29662
rect 8990 29586 9042 29598
rect 10894 29650 10946 29662
rect 10894 29586 10946 29598
rect 11678 29650 11730 29662
rect 11678 29586 11730 29598
rect 14142 29650 14194 29662
rect 14142 29586 14194 29598
rect 17054 29650 17106 29662
rect 17054 29586 17106 29598
rect 17614 29650 17666 29662
rect 17614 29586 17666 29598
rect 19182 29650 19234 29662
rect 19182 29586 19234 29598
rect 20414 29650 20466 29662
rect 20414 29586 20466 29598
rect 24894 29650 24946 29662
rect 24894 29586 24946 29598
rect 25678 29650 25730 29662
rect 25678 29586 25730 29598
rect 34414 29650 34466 29662
rect 57698 29598 57710 29650
rect 57762 29598 57774 29650
rect 34414 29586 34466 29598
rect 12238 29538 12290 29550
rect 19518 29538 19570 29550
rect 18274 29486 18286 29538
rect 18338 29486 18350 29538
rect 12238 29474 12290 29486
rect 19518 29474 19570 29486
rect 26238 29538 26290 29550
rect 26238 29474 26290 29486
rect 10558 29426 10610 29438
rect 10558 29362 10610 29374
rect 10782 29426 10834 29438
rect 10782 29362 10834 29374
rect 11230 29426 11282 29438
rect 11230 29362 11282 29374
rect 18510 29426 18562 29438
rect 18510 29362 18562 29374
rect 18958 29426 19010 29438
rect 18958 29362 19010 29374
rect 22654 29426 22706 29438
rect 22654 29362 22706 29374
rect 23102 29426 23154 29438
rect 23102 29362 23154 29374
rect 23326 29426 23378 29438
rect 58046 29426 58098 29438
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 23326 29362 23378 29374
rect 58046 29362 58098 29374
rect 18174 29314 18226 29326
rect 18174 29250 18226 29262
rect 22206 29314 22258 29326
rect 22206 29250 22258 29262
rect 23214 29314 23266 29326
rect 23214 29250 23266 29262
rect 23774 29314 23826 29326
rect 23774 29250 23826 29262
rect 24222 29314 24274 29326
rect 24222 29250 24274 29262
rect 32174 29314 32226 29326
rect 32174 29250 32226 29262
rect 32734 29314 32786 29326
rect 33730 29262 33742 29314
rect 33794 29262 33806 29314
rect 32734 29250 32786 29262
rect 32846 29202 32898 29214
rect 32846 29138 32898 29150
rect 33966 29202 34018 29214
rect 34178 29150 34190 29202
rect 34242 29199 34254 29202
rect 34402 29199 34414 29202
rect 34242 29153 34414 29199
rect 34242 29150 34254 29153
rect 34402 29150 34414 29153
rect 34466 29150 34478 29202
rect 33966 29138 34018 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 12014 28866 12066 28878
rect 11330 28814 11342 28866
rect 11394 28863 11406 28866
rect 11554 28863 11566 28866
rect 11394 28817 11566 28863
rect 11394 28814 11406 28817
rect 11554 28814 11566 28817
rect 11618 28814 11630 28866
rect 12014 28802 12066 28814
rect 12350 28866 12402 28878
rect 12350 28802 12402 28814
rect 16606 28866 16658 28878
rect 34178 28814 34190 28866
rect 34242 28863 34254 28866
rect 34514 28863 34526 28866
rect 34242 28817 34526 28863
rect 34242 28814 34254 28817
rect 34514 28814 34526 28817
rect 34578 28814 34590 28866
rect 16606 28802 16658 28814
rect 11342 28754 11394 28766
rect 11342 28690 11394 28702
rect 12574 28754 12626 28766
rect 12574 28690 12626 28702
rect 13582 28754 13634 28766
rect 13582 28690 13634 28702
rect 15822 28754 15874 28766
rect 15822 28690 15874 28702
rect 16382 28754 16434 28766
rect 17726 28754 17778 28766
rect 16930 28702 16942 28754
rect 16994 28702 17006 28754
rect 16382 28690 16434 28702
rect 17726 28690 17778 28702
rect 19406 28754 19458 28766
rect 26462 28754 26514 28766
rect 28478 28754 28530 28766
rect 23538 28702 23550 28754
rect 23602 28702 23614 28754
rect 27906 28702 27918 28754
rect 27970 28702 27982 28754
rect 19406 28690 19458 28702
rect 26462 28690 26514 28702
rect 28478 28690 28530 28702
rect 33294 28754 33346 28766
rect 33294 28690 33346 28702
rect 34190 28754 34242 28766
rect 34190 28690 34242 28702
rect 34638 28754 34690 28766
rect 34638 28690 34690 28702
rect 35758 28754 35810 28766
rect 35758 28690 35810 28702
rect 58158 28754 58210 28766
rect 58158 28690 58210 28702
rect 18174 28642 18226 28654
rect 18174 28578 18226 28590
rect 18286 28642 18338 28654
rect 18286 28578 18338 28590
rect 18734 28642 18786 28654
rect 18734 28578 18786 28590
rect 18958 28642 19010 28654
rect 24222 28642 24274 28654
rect 23090 28590 23102 28642
rect 23154 28590 23166 28642
rect 23426 28590 23438 28642
rect 23490 28590 23502 28642
rect 18958 28578 19010 28590
rect 24222 28578 24274 28590
rect 24670 28642 24722 28654
rect 35982 28642 36034 28654
rect 27458 28590 27470 28642
rect 27522 28590 27534 28642
rect 24670 28578 24722 28590
rect 35982 28578 36034 28590
rect 38110 28642 38162 28654
rect 38110 28578 38162 28590
rect 38558 28642 38610 28654
rect 38558 28578 38610 28590
rect 39566 28642 39618 28654
rect 40462 28642 40514 28654
rect 39890 28590 39902 28642
rect 39954 28590 39966 28642
rect 39566 28578 39618 28590
rect 40462 28578 40514 28590
rect 42254 28642 42306 28654
rect 42254 28578 42306 28590
rect 18510 28530 18562 28542
rect 18510 28466 18562 28478
rect 27022 28530 27074 28542
rect 27022 28466 27074 28478
rect 35310 28530 35362 28542
rect 35310 28466 35362 28478
rect 35534 28530 35586 28542
rect 35534 28466 35586 28478
rect 39118 28530 39170 28542
rect 39330 28478 39342 28530
rect 39394 28478 39406 28530
rect 41346 28478 41358 28530
rect 41410 28478 41422 28530
rect 39118 28466 39170 28478
rect 35422 28418 35474 28430
rect 22978 28366 22990 28418
rect 23042 28366 23054 28418
rect 35422 28354 35474 28366
rect 39902 28418 39954 28430
rect 39902 28354 39954 28366
rect 41694 28418 41746 28430
rect 41694 28354 41746 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 6078 28082 6130 28094
rect 6078 28018 6130 28030
rect 7310 28082 7362 28094
rect 7310 28018 7362 28030
rect 10894 28082 10946 28094
rect 10894 28018 10946 28030
rect 12014 28082 12066 28094
rect 12014 28018 12066 28030
rect 12910 28082 12962 28094
rect 12910 28018 12962 28030
rect 17726 28082 17778 28094
rect 17726 28018 17778 28030
rect 23326 28082 23378 28094
rect 23326 28018 23378 28030
rect 28702 28082 28754 28094
rect 28702 28018 28754 28030
rect 29262 28082 29314 28094
rect 29262 28018 29314 28030
rect 23214 27970 23266 27982
rect 23214 27906 23266 27918
rect 23774 27970 23826 27982
rect 23774 27906 23826 27918
rect 24222 27970 24274 27982
rect 24222 27906 24274 27918
rect 28814 27970 28866 27982
rect 28814 27906 28866 27918
rect 6302 27858 6354 27870
rect 6302 27794 6354 27806
rect 6750 27858 6802 27870
rect 6750 27794 6802 27806
rect 10558 27858 10610 27870
rect 10558 27794 10610 27806
rect 10782 27858 10834 27870
rect 10782 27794 10834 27806
rect 11006 27858 11058 27870
rect 11006 27794 11058 27806
rect 11566 27858 11618 27870
rect 11566 27794 11618 27806
rect 23550 27858 23602 27870
rect 23550 27794 23602 27806
rect 10110 27746 10162 27758
rect 6066 27694 6078 27746
rect 6130 27694 6142 27746
rect 10110 27682 10162 27694
rect 24670 27746 24722 27758
rect 24670 27682 24722 27694
rect 10334 27634 10386 27646
rect 10334 27570 10386 27582
rect 28702 27634 28754 27646
rect 28702 27570 28754 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 18734 27298 18786 27310
rect 18734 27234 18786 27246
rect 25342 27298 25394 27310
rect 25342 27234 25394 27246
rect 34078 27298 34130 27310
rect 34078 27234 34130 27246
rect 3502 27186 3554 27198
rect 3502 27122 3554 27134
rect 11454 27186 11506 27198
rect 11454 27122 11506 27134
rect 17838 27186 17890 27198
rect 17838 27122 17890 27134
rect 18286 27186 18338 27198
rect 18286 27122 18338 27134
rect 20190 27186 20242 27198
rect 26014 27186 26066 27198
rect 24546 27134 24558 27186
rect 24610 27134 24622 27186
rect 20190 27122 20242 27134
rect 26014 27122 26066 27134
rect 29486 27186 29538 27198
rect 29486 27122 29538 27134
rect 31278 27186 31330 27198
rect 31278 27122 31330 27134
rect 12126 27074 12178 27086
rect 3042 27022 3054 27074
rect 3106 27022 3118 27074
rect 11666 27022 11678 27074
rect 11730 27022 11742 27074
rect 12126 27010 12178 27022
rect 17390 27074 17442 27086
rect 19406 27074 19458 27086
rect 19170 27022 19182 27074
rect 19234 27022 19246 27074
rect 17390 27010 17442 27022
rect 19406 27010 19458 27022
rect 19630 27074 19682 27086
rect 19630 27010 19682 27022
rect 22878 27074 22930 27086
rect 22878 27010 22930 27022
rect 23326 27074 23378 27086
rect 23326 27010 23378 27022
rect 23550 27074 23602 27086
rect 23550 27010 23602 27022
rect 24446 27074 24498 27086
rect 25118 27074 25170 27086
rect 31726 27074 31778 27086
rect 24770 27022 24782 27074
rect 24834 27022 24846 27074
rect 27682 27022 27694 27074
rect 27746 27022 27758 27074
rect 28018 27022 28030 27074
rect 28082 27022 28094 27074
rect 32722 27022 32734 27074
rect 32786 27022 32798 27074
rect 33282 27022 33294 27074
rect 33346 27022 33358 27074
rect 33730 27022 33742 27074
rect 33794 27022 33806 27074
rect 24446 27010 24498 27022
rect 25118 27010 25170 27022
rect 31726 27010 31778 27022
rect 11342 26962 11394 26974
rect 2146 26910 2158 26962
rect 2210 26910 2222 26962
rect 11342 26898 11394 26910
rect 19518 26962 19570 26974
rect 19518 26898 19570 26910
rect 24670 26962 24722 26974
rect 24670 26898 24722 26910
rect 26462 26962 26514 26974
rect 27010 26910 27022 26962
rect 27074 26910 27086 26962
rect 28578 26910 28590 26962
rect 28642 26910 28654 26962
rect 32610 26910 32622 26962
rect 32674 26910 32686 26962
rect 26462 26898 26514 26910
rect 23214 26850 23266 26862
rect 28466 26798 28478 26850
rect 28530 26798 28542 26850
rect 23214 26786 23266 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 10222 26514 10274 26526
rect 10222 26450 10274 26462
rect 11342 26514 11394 26526
rect 11342 26450 11394 26462
rect 12462 26514 12514 26526
rect 12462 26450 12514 26462
rect 23662 26514 23714 26526
rect 23662 26450 23714 26462
rect 23998 26514 24050 26526
rect 23998 26450 24050 26462
rect 24558 26514 24610 26526
rect 24558 26450 24610 26462
rect 25678 26514 25730 26526
rect 25678 26450 25730 26462
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 27806 26514 27858 26526
rect 27806 26450 27858 26462
rect 32174 26514 32226 26526
rect 32174 26450 32226 26462
rect 42030 26514 42082 26526
rect 42030 26450 42082 26462
rect 42702 26514 42754 26526
rect 42702 26450 42754 26462
rect 12014 26402 12066 26414
rect 12014 26338 12066 26350
rect 27022 26402 27074 26414
rect 27022 26338 27074 26350
rect 41582 26402 41634 26414
rect 41582 26338 41634 26350
rect 10782 26290 10834 26302
rect 10782 26226 10834 26238
rect 41918 26290 41970 26302
rect 41918 26226 41970 26238
rect 42142 26290 42194 26302
rect 42142 26226 42194 26238
rect 43038 26178 43090 26190
rect 27346 26126 27358 26178
rect 27410 26126 27422 26178
rect 43038 26114 43090 26126
rect 11902 26066 11954 26078
rect 42354 26014 42366 26066
rect 42418 26063 42430 26066
rect 43026 26063 43038 26066
rect 42418 26017 43038 26063
rect 42418 26014 42430 26017
rect 43026 26014 43038 26017
rect 43090 26014 43102 26066
rect 11902 26002 11954 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 22542 25730 22594 25742
rect 22542 25666 22594 25678
rect 24110 25730 24162 25742
rect 24110 25666 24162 25678
rect 11566 25618 11618 25630
rect 9762 25566 9774 25618
rect 9826 25566 9838 25618
rect 10658 25566 10670 25618
rect 10722 25566 10734 25618
rect 11566 25554 11618 25566
rect 22430 25618 22482 25630
rect 22430 25554 22482 25566
rect 22990 25618 23042 25630
rect 22990 25554 23042 25566
rect 56254 25618 56306 25630
rect 57810 25566 57822 25618
rect 57874 25566 57886 25618
rect 56254 25554 56306 25566
rect 10882 25454 10894 25506
rect 10946 25454 10958 25506
rect 56802 25454 56814 25506
rect 56866 25454 56878 25506
rect 9774 25394 9826 25406
rect 9774 25330 9826 25342
rect 9998 25394 10050 25406
rect 9998 25330 10050 25342
rect 23998 25394 24050 25406
rect 23998 25330 24050 25342
rect 24110 25282 24162 25294
rect 24110 25218 24162 25230
rect 24670 25282 24722 25294
rect 24670 25218 24722 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 9774 24946 9826 24958
rect 9774 24882 9826 24894
rect 10334 24946 10386 24958
rect 10334 24882 10386 24894
rect 10782 24946 10834 24958
rect 10782 24882 10834 24894
rect 19742 24946 19794 24958
rect 19742 24882 19794 24894
rect 21758 24946 21810 24958
rect 21758 24882 21810 24894
rect 22318 24946 22370 24958
rect 22318 24882 22370 24894
rect 23214 24946 23266 24958
rect 23214 24882 23266 24894
rect 24670 24946 24722 24958
rect 24670 24882 24722 24894
rect 24782 24946 24834 24958
rect 24782 24882 24834 24894
rect 26910 24946 26962 24958
rect 26910 24882 26962 24894
rect 27470 24946 27522 24958
rect 27470 24882 27522 24894
rect 27806 24946 27858 24958
rect 27806 24882 27858 24894
rect 28254 24946 28306 24958
rect 28254 24882 28306 24894
rect 28366 24946 28418 24958
rect 28366 24882 28418 24894
rect 28590 24946 28642 24958
rect 28590 24882 28642 24894
rect 10894 24834 10946 24846
rect 10894 24770 10946 24782
rect 11342 24834 11394 24846
rect 11342 24770 11394 24782
rect 12238 24834 12290 24846
rect 12238 24770 12290 24782
rect 28814 24834 28866 24846
rect 28814 24770 28866 24782
rect 11106 24670 11118 24722
rect 11170 24670 11182 24722
rect 24210 24670 24222 24722
rect 24274 24670 24286 24722
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 11790 24610 11842 24622
rect 11790 24546 11842 24558
rect 19630 24610 19682 24622
rect 19630 24546 19682 24558
rect 22430 24610 22482 24622
rect 22430 24546 22482 24558
rect 23662 24610 23714 24622
rect 23662 24546 23714 24558
rect 9762 24446 9774 24498
rect 9826 24495 9838 24498
rect 10658 24495 10670 24498
rect 9826 24449 10670 24495
rect 9826 24446 9838 24449
rect 10658 24446 10670 24449
rect 10722 24446 10734 24498
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 3614 24050 3666 24062
rect 3614 23986 3666 23998
rect 18174 24050 18226 24062
rect 18174 23986 18226 23998
rect 18622 24050 18674 24062
rect 26350 24050 26402 24062
rect 25106 23998 25118 24050
rect 25170 23998 25182 24050
rect 18622 23986 18674 23998
rect 26350 23986 26402 23998
rect 17166 23938 17218 23950
rect 3042 23886 3054 23938
rect 3106 23886 3118 23938
rect 17166 23874 17218 23886
rect 17390 23938 17442 23950
rect 22754 23886 22766 23938
rect 22818 23886 22830 23938
rect 24322 23886 24334 23938
rect 24386 23886 24398 23938
rect 17390 23874 17442 23886
rect 2146 23774 2158 23826
rect 2210 23774 2222 23826
rect 17714 23774 17726 23826
rect 17778 23774 17790 23826
rect 23202 23774 23214 23826
rect 23266 23774 23278 23826
rect 24210 23774 24222 23826
rect 24274 23774 24286 23826
rect 21646 23714 21698 23726
rect 21646 23650 21698 23662
rect 22094 23714 22146 23726
rect 22094 23650 22146 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 11342 23378 11394 23390
rect 11342 23314 11394 23326
rect 18062 23378 18114 23390
rect 18062 23314 18114 23326
rect 18846 23378 18898 23390
rect 18846 23314 18898 23326
rect 19182 23378 19234 23390
rect 19182 23314 19234 23326
rect 21198 23378 21250 23390
rect 21198 23314 21250 23326
rect 22094 23378 22146 23390
rect 22094 23314 22146 23326
rect 23550 23378 23602 23390
rect 23550 23314 23602 23326
rect 9774 23266 9826 23278
rect 9774 23202 9826 23214
rect 17950 23266 18002 23278
rect 57710 23266 57762 23278
rect 22978 23214 22990 23266
rect 23042 23214 23054 23266
rect 17950 23202 18002 23214
rect 57710 23202 57762 23214
rect 17838 23154 17890 23166
rect 10434 23102 10446 23154
rect 10498 23102 10510 23154
rect 17838 23090 17890 23102
rect 18398 23154 18450 23166
rect 18398 23090 18450 23102
rect 22318 23154 22370 23166
rect 22318 23090 22370 23102
rect 22766 23154 22818 23166
rect 22766 23090 22818 23102
rect 23102 23154 23154 23166
rect 23102 23090 23154 23102
rect 58046 23154 58098 23166
rect 58046 23090 58098 23102
rect 11678 23042 11730 23054
rect 10658 22990 10670 23042
rect 10722 22990 10734 23042
rect 11678 22978 11730 22990
rect 16942 23042 16994 23054
rect 16942 22978 16994 22990
rect 21646 23042 21698 23054
rect 21646 22978 21698 22990
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 10994 22542 11006 22594
rect 11058 22542 11070 22594
rect 9438 22482 9490 22494
rect 9438 22418 9490 22430
rect 11790 22482 11842 22494
rect 11790 22418 11842 22430
rect 58158 22482 58210 22494
rect 58158 22418 58210 22430
rect 10110 22370 10162 22382
rect 10110 22306 10162 22318
rect 10334 22370 10386 22382
rect 10334 22306 10386 22318
rect 10558 22370 10610 22382
rect 10558 22306 10610 22318
rect 12238 22370 12290 22382
rect 12238 22306 12290 22318
rect 9998 22258 10050 22270
rect 9998 22194 10050 22206
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 3502 21810 3554 21822
rect 3502 21746 3554 21758
rect 11342 21810 11394 21822
rect 11342 21746 11394 21758
rect 3042 21534 3054 21586
rect 3106 21534 3118 21586
rect 2034 21422 2046 21474
rect 2098 21422 2110 21474
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 4286 20914 4338 20926
rect 4286 20850 4338 20862
rect 57710 20690 57762 20702
rect 57710 20626 57762 20638
rect 58046 20690 58098 20702
rect 58046 20626 58098 20638
rect 3726 20578 3778 20590
rect 3726 20514 3778 20526
rect 57262 20578 57314 20590
rect 57262 20514 57314 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 1822 17554 1874 17566
rect 1822 17490 1874 17502
rect 2158 17554 2210 17566
rect 2158 17490 2210 17502
rect 57710 17554 57762 17566
rect 57710 17490 57762 17502
rect 58046 17554 58098 17566
rect 58046 17490 58098 17502
rect 57262 17442 57314 17454
rect 57262 17378 57314 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 1822 17106 1874 17118
rect 1822 17042 1874 17054
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 2158 15538 2210 15550
rect 2158 15474 2210 15486
rect 1822 15314 1874 15326
rect 1822 15250 1874 15262
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 1822 14642 1874 14654
rect 1822 14578 1874 14590
rect 56366 14642 56418 14654
rect 56366 14578 56418 14590
rect 56802 14478 56814 14530
rect 56866 14478 56878 14530
rect 57698 14366 57710 14418
rect 57762 14366 57774 14418
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 3502 12402 3554 12414
rect 3502 12338 3554 12350
rect 3042 12126 3054 12178
rect 3106 12126 3118 12178
rect 2034 12014 2046 12066
rect 2098 12014 2110 12066
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 56802 11342 56814 11394
rect 56866 11342 56878 11394
rect 57698 11230 57710 11282
rect 57762 11230 57774 11282
rect 56366 11170 56418 11182
rect 56366 11106 56418 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 2158 9266 2210 9278
rect 2158 9202 2210 9214
rect 1822 9042 1874 9054
rect 1822 8978 1874 8990
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 1822 8370 1874 8382
rect 1822 8306 1874 8318
rect 57710 8146 57762 8158
rect 57710 8082 57762 8094
rect 58046 8146 58098 8158
rect 58046 8082 58098 8094
rect 57262 8034 57314 8046
rect 57262 7970 57314 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 3502 6130 3554 6142
rect 3502 6066 3554 6078
rect 58046 6018 58098 6030
rect 58046 5954 58098 5966
rect 3042 5854 3054 5906
rect 3106 5854 3118 5906
rect 2034 5742 2046 5794
rect 2098 5742 2110 5794
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 3614 5234 3666 5246
rect 3614 5170 3666 5182
rect 3042 5070 3054 5122
rect 3106 5070 3118 5122
rect 57262 5010 57314 5022
rect 2146 4958 2158 5010
rect 2210 4958 2222 5010
rect 57262 4946 57314 4958
rect 57710 5010 57762 5022
rect 57710 4946 57762 4958
rect 58046 5010 58098 5022
rect 58046 4946 58098 4958
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 3502 4562 3554 4574
rect 3502 4498 3554 4510
rect 4398 4562 4450 4574
rect 4398 4498 4450 4510
rect 11118 4562 11170 4574
rect 11118 4498 11170 4510
rect 16494 4562 16546 4574
rect 16494 4498 16546 4510
rect 34750 4562 34802 4574
rect 34750 4498 34802 4510
rect 57710 4562 57762 4574
rect 57710 4498 57762 4510
rect 58046 4338 58098 4350
rect 3042 4286 3054 4338
rect 3106 4286 3118 4338
rect 58046 4274 58098 4286
rect 56814 4226 56866 4238
rect 2034 4174 2046 4226
rect 2098 4174 2110 4226
rect 56814 4162 56866 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 16830 3666 16882 3678
rect 32510 3666 32562 3678
rect 44270 3666 44322 3678
rect 15250 3614 15262 3666
rect 15314 3614 15326 3666
rect 18386 3614 18398 3666
rect 18450 3614 18462 3666
rect 35746 3614 35758 3666
rect 35810 3614 35822 3666
rect 45154 3614 45166 3666
rect 45218 3614 45230 3666
rect 16830 3602 16882 3614
rect 32510 3602 32562 3614
rect 44270 3602 44322 3614
rect 56030 3554 56082 3566
rect 4162 3502 4174 3554
rect 4226 3502 4238 3554
rect 10882 3502 10894 3554
rect 10946 3502 10958 3554
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 17714 3502 17726 3554
rect 17778 3502 17790 3554
rect 33170 3502 33182 3554
rect 33234 3502 33246 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 45938 3502 45950 3554
rect 46002 3502 46014 3554
rect 56690 3502 56702 3554
rect 56754 3502 56766 3554
rect 56030 3490 56082 3502
rect 5070 3442 5122 3454
rect 3266 3390 3278 3442
rect 3330 3390 3342 3442
rect 5070 3378 5122 3390
rect 5742 3442 5794 3454
rect 20750 3442 20802 3454
rect 9986 3390 9998 3442
rect 10050 3390 10062 3442
rect 5742 3378 5794 3390
rect 20750 3378 20802 3390
rect 21422 3442 21474 3454
rect 21422 3378 21474 3390
rect 23326 3442 23378 3454
rect 23326 3378 23378 3390
rect 23774 3442 23826 3454
rect 23774 3378 23826 3390
rect 29374 3442 29426 3454
rect 29374 3378 29426 3390
rect 29822 3442 29874 3454
rect 41470 3442 41522 3454
rect 34066 3390 34078 3442
rect 34130 3390 34142 3442
rect 29822 3378 29874 3390
rect 41470 3378 41522 3390
rect 41918 3442 41970 3454
rect 41918 3378 41970 3390
rect 48190 3442 48242 3454
rect 48190 3378 48242 3390
rect 49198 3442 49250 3454
rect 49198 3378 49250 3390
rect 50206 3442 50258 3454
rect 50206 3378 50258 3390
rect 50990 3442 51042 3454
rect 57586 3390 57598 3442
rect 57650 3390 57662 3442
rect 50990 3378 51042 3390
rect 6078 3330 6130 3342
rect 6078 3266 6130 3278
rect 11678 3330 11730 3342
rect 11678 3266 11730 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 24110 3330 24162 3342
rect 24110 3266 24162 3278
rect 27134 3330 27186 3342
rect 27134 3266 27186 3278
rect 30158 3330 30210 3342
rect 30158 3266 30210 3278
rect 42254 3330 42306 3342
rect 42254 3266 42306 3278
rect 48862 3330 48914 3342
rect 48862 3266 48914 3278
rect 50654 3330 50706 3342
rect 50654 3266 50706 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 29038 56590 29090 56642
rect 29934 56590 29986 56642
rect 52334 56590 52386 56642
rect 53006 56590 53058 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 8318 56254 8370 56306
rect 19294 56254 19346 56306
rect 31390 56254 31442 56306
rect 34750 56254 34802 56306
rect 37438 56254 37490 56306
rect 46174 56254 46226 56306
rect 52110 56254 52162 56306
rect 55134 56254 55186 56306
rect 2606 56142 2658 56194
rect 6078 56142 6130 56194
rect 11342 56142 11394 56194
rect 19742 56142 19794 56194
rect 20078 56142 20130 56194
rect 23438 56142 23490 56194
rect 26126 56142 26178 56194
rect 31838 56142 31890 56194
rect 35198 56142 35250 56194
rect 35534 56142 35586 56194
rect 37886 56142 37938 56194
rect 38222 56142 38274 56194
rect 42142 56142 42194 56194
rect 46622 56142 46674 56194
rect 52782 56142 52834 56194
rect 55582 56142 55634 56194
rect 55918 56142 55970 56194
rect 57710 56142 57762 56194
rect 3502 56030 3554 56082
rect 6974 56030 7026 56082
rect 7534 56030 7586 56082
rect 12238 56030 12290 56082
rect 18734 56030 18786 56082
rect 24110 56030 24162 56082
rect 25342 56030 25394 56082
rect 26798 56030 26850 56082
rect 29262 56030 29314 56082
rect 32062 56030 32114 56082
rect 41246 56030 41298 56082
rect 46846 56030 46898 56082
rect 49534 56030 49586 56082
rect 49982 56030 50034 56082
rect 53006 56030 53058 56082
rect 56814 56030 56866 56082
rect 4062 55918 4114 55970
rect 12798 55918 12850 55970
rect 17726 55918 17778 55970
rect 20638 55918 20690 55970
rect 22654 55918 22706 55970
rect 28590 55918 28642 55970
rect 29934 55918 29986 55970
rect 40350 55918 40402 55970
rect 50654 55918 50706 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 55806 55470 55858 55522
rect 56590 55470 56642 55522
rect 57822 55358 57874 55410
rect 10782 55246 10834 55298
rect 11342 55246 11394 55298
rect 15822 55246 15874 55298
rect 16270 55246 16322 55298
rect 56814 55246 56866 55298
rect 1822 55134 1874 55186
rect 2158 55022 2210 55074
rect 7646 55022 7698 55074
rect 8318 55022 8370 55074
rect 11902 55022 11954 55074
rect 12350 55022 12402 55074
rect 18734 55022 18786 55074
rect 19294 55022 19346 55074
rect 19854 55022 19906 55074
rect 20302 55022 20354 55074
rect 20862 55022 20914 55074
rect 55806 55022 55858 55074
rect 56254 55022 56306 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 1822 54686 1874 54738
rect 23214 54686 23266 54738
rect 58046 54686 58098 54738
rect 20078 54462 20130 54514
rect 20750 54462 20802 54514
rect 11454 54350 11506 54402
rect 12350 54350 12402 54402
rect 19630 54350 19682 54402
rect 24222 54350 24274 54402
rect 27806 54350 27858 54402
rect 29150 54350 29202 54402
rect 30718 54350 30770 54402
rect 23774 54238 23826 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 30270 53902 30322 53954
rect 38894 53902 38946 53954
rect 39790 53902 39842 53954
rect 3726 53790 3778 53842
rect 27470 53790 27522 53842
rect 39230 53790 39282 53842
rect 42366 53790 42418 53842
rect 4062 53678 4114 53730
rect 4622 53678 4674 53730
rect 8654 53678 8706 53730
rect 9102 53678 9154 53730
rect 14478 53678 14530 53730
rect 14814 53678 14866 53730
rect 18734 53678 18786 53730
rect 28702 53678 28754 53730
rect 32510 53678 32562 53730
rect 32622 53678 32674 53730
rect 33070 53678 33122 53730
rect 38446 53678 38498 53730
rect 41582 53678 41634 53730
rect 41918 53678 41970 53730
rect 42142 53678 42194 53730
rect 1822 53566 1874 53618
rect 12126 53566 12178 53618
rect 27358 53566 27410 53618
rect 28814 53566 28866 53618
rect 30382 53566 30434 53618
rect 31054 53566 31106 53618
rect 42814 53566 42866 53618
rect 45614 53566 45666 53618
rect 2158 53454 2210 53506
rect 3838 53454 3890 53506
rect 11566 53454 11618 53506
rect 12686 53454 12738 53506
rect 13806 53454 13858 53506
rect 17390 53454 17442 53506
rect 17950 53454 18002 53506
rect 18286 53454 18338 53506
rect 28254 53454 28306 53506
rect 29486 53454 29538 53506
rect 30942 53454 30994 53506
rect 31502 53454 31554 53506
rect 39118 53454 39170 53506
rect 39902 53454 39954 53506
rect 40014 53454 40066 53506
rect 40686 53454 40738 53506
rect 41470 53454 41522 53506
rect 41694 53454 41746 53506
rect 45502 53454 45554 53506
rect 46062 53454 46114 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 1822 53118 1874 53170
rect 23438 53118 23490 53170
rect 29038 53118 29090 53170
rect 29710 53118 29762 53170
rect 3726 53006 3778 53058
rect 3950 53006 4002 53058
rect 6190 53006 6242 53058
rect 14142 53006 14194 53058
rect 18622 53006 18674 53058
rect 28030 53006 28082 53058
rect 28254 53006 28306 53058
rect 30494 53006 30546 53058
rect 31166 53006 31218 53058
rect 42702 53006 42754 53058
rect 43374 53006 43426 53058
rect 8542 52894 8594 52946
rect 9102 52894 9154 52946
rect 16494 52894 16546 52946
rect 17054 52894 17106 52946
rect 20526 52894 20578 52946
rect 21086 52894 21138 52946
rect 31614 52894 31666 52946
rect 3838 52782 3890 52834
rect 4510 52782 4562 52834
rect 9662 52782 9714 52834
rect 10222 52782 10274 52834
rect 10558 52782 10610 52834
rect 12462 52782 12514 52834
rect 17614 52782 17666 52834
rect 18174 52782 18226 52834
rect 19966 52782 20018 52834
rect 24558 52782 24610 52834
rect 27358 52782 27410 52834
rect 29150 52782 29202 52834
rect 29822 52782 29874 52834
rect 39454 52782 39506 52834
rect 40798 52782 40850 52834
rect 41470 52782 41522 52834
rect 43598 52782 43650 52834
rect 44046 52782 44098 52834
rect 5406 52670 5458 52722
rect 13358 52670 13410 52722
rect 24110 52670 24162 52722
rect 27246 52670 27298 52722
rect 27918 52670 27970 52722
rect 30382 52670 30434 52722
rect 31054 52670 31106 52722
rect 43262 52670 43314 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 31390 52334 31442 52386
rect 51438 52334 51490 52386
rect 11902 52222 11954 52274
rect 20526 52222 20578 52274
rect 21534 52222 21586 52274
rect 28478 52222 28530 52274
rect 29486 52222 29538 52274
rect 30046 52222 30098 52274
rect 30718 52222 30770 52274
rect 31502 52222 31554 52274
rect 52670 52222 52722 52274
rect 7198 52110 7250 52162
rect 10222 52110 10274 52162
rect 10894 52110 10946 52162
rect 11454 52110 11506 52162
rect 16494 52110 16546 52162
rect 16942 52110 16994 52162
rect 22094 52110 22146 52162
rect 27582 52110 27634 52162
rect 28366 52110 28418 52162
rect 51774 52110 51826 52162
rect 52222 52110 52274 52162
rect 53454 52110 53506 52162
rect 53566 52110 53618 52162
rect 54126 52110 54178 52162
rect 7982 51886 8034 51938
rect 19182 51886 19234 51938
rect 19966 51886 20018 51938
rect 31950 51886 32002 51938
rect 51550 51886 51602 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 22654 51550 22706 51602
rect 40126 51550 40178 51602
rect 53118 51550 53170 51602
rect 3950 51438 4002 51490
rect 4622 51438 4674 51490
rect 18734 51438 18786 51490
rect 11118 51326 11170 51378
rect 19518 51326 19570 51378
rect 20190 51326 20242 51378
rect 39902 51326 39954 51378
rect 40238 51326 40290 51378
rect 40798 51326 40850 51378
rect 43150 51326 43202 51378
rect 43486 51326 43538 51378
rect 5182 51214 5234 51266
rect 11902 51214 11954 51266
rect 18286 51214 18338 51266
rect 23662 51214 23714 51266
rect 38558 51214 38610 51266
rect 39006 51214 39058 51266
rect 40014 51214 40066 51266
rect 41582 51214 41634 51266
rect 42142 51214 42194 51266
rect 42478 51214 42530 51266
rect 43038 51214 43090 51266
rect 3726 51102 3778 51154
rect 4062 51102 4114 51154
rect 4734 51102 4786 51154
rect 23214 51102 23266 51154
rect 40574 51102 40626 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 39118 50766 39170 50818
rect 39790 50766 39842 50818
rect 40462 50766 40514 50818
rect 18622 50654 18674 50706
rect 35534 50654 35586 50706
rect 40126 50654 40178 50706
rect 8206 50542 8258 50594
rect 8654 50542 8706 50594
rect 15038 50542 15090 50594
rect 15598 50542 15650 50594
rect 19742 50542 19794 50594
rect 1822 50430 1874 50482
rect 12238 50430 12290 50482
rect 12686 50430 12738 50482
rect 39454 50430 39506 50482
rect 40238 50430 40290 50482
rect 40910 50430 40962 50482
rect 57262 50430 57314 50482
rect 58046 50430 58098 50482
rect 2158 50318 2210 50370
rect 11118 50318 11170 50370
rect 11678 50318 11730 50370
rect 18062 50318 18114 50370
rect 19182 50318 19234 50370
rect 32398 50318 32450 50370
rect 36094 50318 36146 50370
rect 36654 50318 36706 50370
rect 57710 50318 57762 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 1822 49982 1874 50034
rect 22094 49982 22146 50034
rect 43598 49982 43650 50034
rect 44270 49982 44322 50034
rect 44942 49982 44994 50034
rect 12238 49870 12290 49922
rect 32174 49870 32226 49922
rect 32622 49870 32674 49922
rect 35870 49870 35922 49922
rect 44494 49870 44546 49922
rect 15038 49758 15090 49810
rect 18958 49758 19010 49810
rect 19630 49758 19682 49810
rect 36430 49758 36482 49810
rect 15598 49646 15650 49698
rect 18510 49646 18562 49698
rect 23102 49646 23154 49698
rect 31502 49646 31554 49698
rect 36878 49646 36930 49698
rect 22654 49534 22706 49586
rect 31390 49534 31442 49586
rect 32062 49534 32114 49586
rect 44158 49534 44210 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 27694 49198 27746 49250
rect 27918 49198 27970 49250
rect 11006 49086 11058 49138
rect 18510 49086 18562 49138
rect 27918 49086 27970 49138
rect 31950 49086 32002 49138
rect 32398 49086 32450 49138
rect 35870 49086 35922 49138
rect 9774 48974 9826 49026
rect 10334 48974 10386 49026
rect 20526 48974 20578 49026
rect 31838 48862 31890 48914
rect 6638 48750 6690 48802
rect 7422 48750 7474 48802
rect 11342 48750 11394 48802
rect 21534 48750 21586 48802
rect 36430 48750 36482 48802
rect 37438 48750 37490 48802
rect 47518 48750 47570 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4510 48414 4562 48466
rect 10558 48414 10610 48466
rect 12126 48414 12178 48466
rect 46622 48414 46674 48466
rect 47070 48414 47122 48466
rect 3950 48302 4002 48354
rect 27694 48302 27746 48354
rect 48078 48302 48130 48354
rect 48190 48302 48242 48354
rect 3054 48190 3106 48242
rect 37998 48190 38050 48242
rect 47854 48190 47906 48242
rect 2046 48078 2098 48130
rect 3950 48078 4002 48130
rect 28702 48078 28754 48130
rect 29150 48078 29202 48130
rect 38558 48078 38610 48130
rect 3726 47966 3778 48018
rect 27582 47966 27634 48018
rect 28590 47966 28642 48018
rect 37886 47966 37938 48018
rect 48638 47966 48690 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 18398 47518 18450 47570
rect 19406 47518 19458 47570
rect 26798 47518 26850 47570
rect 27358 47518 27410 47570
rect 46846 47518 46898 47570
rect 47294 47518 47346 47570
rect 49086 47518 49138 47570
rect 8542 47406 8594 47458
rect 8990 47406 9042 47458
rect 14030 47406 14082 47458
rect 28030 47406 28082 47458
rect 48078 47406 48130 47458
rect 48302 47406 48354 47458
rect 48750 47406 48802 47458
rect 28702 47294 28754 47346
rect 3278 47182 3330 47234
rect 11454 47182 11506 47234
rect 12014 47182 12066 47234
rect 12574 47182 12626 47234
rect 27246 47182 27298 47234
rect 27918 47182 27970 47234
rect 28590 47182 28642 47234
rect 29486 47182 29538 47234
rect 48414 47182 48466 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4510 46846 4562 46898
rect 23438 46846 23490 46898
rect 28254 46846 28306 46898
rect 28702 46846 28754 46898
rect 29934 46846 29986 46898
rect 43038 46846 43090 46898
rect 4062 46734 4114 46786
rect 27806 46734 27858 46786
rect 29486 46734 29538 46786
rect 3726 46622 3778 46674
rect 20414 46622 20466 46674
rect 21086 46622 21138 46674
rect 42926 46622 42978 46674
rect 43150 46622 43202 46674
rect 43822 46622 43874 46674
rect 47966 46622 48018 46674
rect 3166 46510 3218 46562
rect 9774 46510 9826 46562
rect 12350 46510 12402 46562
rect 19630 46510 19682 46562
rect 20078 46510 20130 46562
rect 24558 46510 24610 46562
rect 29374 46510 29426 46562
rect 32958 46510 33010 46562
rect 33742 46510 33794 46562
rect 34414 46510 34466 46562
rect 34862 46510 34914 46562
rect 37102 46510 37154 46562
rect 37438 46510 37490 46562
rect 41806 46510 41858 46562
rect 42366 46510 42418 46562
rect 43374 46510 43426 46562
rect 47742 46510 47794 46562
rect 48078 46510 48130 46562
rect 48750 46510 48802 46562
rect 3726 46398 3778 46450
rect 24110 46398 24162 46450
rect 27694 46398 27746 46450
rect 33630 46398 33682 46450
rect 34302 46398 34354 46450
rect 43598 46398 43650 46450
rect 47630 46398 47682 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 35870 46062 35922 46114
rect 38334 46062 38386 46114
rect 11230 45950 11282 46002
rect 31726 45950 31778 46002
rect 32398 45950 32450 46002
rect 35422 45950 35474 46002
rect 10110 45838 10162 45890
rect 10670 45838 10722 45890
rect 11678 45838 11730 45890
rect 19182 45838 19234 45890
rect 19630 45838 19682 45890
rect 30718 45838 30770 45890
rect 35534 45838 35586 45890
rect 35758 45838 35810 45890
rect 36206 45838 36258 45890
rect 37998 45838 38050 45890
rect 38558 45838 38610 45890
rect 16158 45726 16210 45778
rect 16942 45726 16994 45778
rect 34078 45726 34130 45778
rect 34526 45726 34578 45778
rect 6974 45614 7026 45666
rect 7758 45614 7810 45666
rect 20414 45614 20466 45666
rect 20862 45614 20914 45666
rect 28702 45614 28754 45666
rect 30606 45614 30658 45666
rect 31166 45614 31218 45666
rect 33966 45614 34018 45666
rect 35982 45614 36034 45666
rect 36654 45614 36706 45666
rect 37662 45614 37714 45666
rect 37774 45614 37826 45666
rect 37886 45614 37938 45666
rect 39006 45614 39058 45666
rect 40350 45614 40402 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2158 45278 2210 45330
rect 23326 45278 23378 45330
rect 27582 45278 27634 45330
rect 29934 45278 29986 45330
rect 30718 45278 30770 45330
rect 32622 45278 32674 45330
rect 39902 45278 39954 45330
rect 40798 45278 40850 45330
rect 6190 45166 6242 45218
rect 31502 45166 31554 45218
rect 32174 45166 32226 45218
rect 37326 45166 37378 45218
rect 38222 45166 38274 45218
rect 39790 45166 39842 45218
rect 40686 45166 40738 45218
rect 1822 45054 1874 45106
rect 8542 45054 8594 45106
rect 8878 45054 8930 45106
rect 11230 45054 11282 45106
rect 20190 45054 20242 45106
rect 20750 45054 20802 45106
rect 29262 45054 29314 45106
rect 29710 45054 29762 45106
rect 30158 45054 30210 45106
rect 36990 45054 37042 45106
rect 9774 44942 9826 44994
rect 10110 44942 10162 44994
rect 10782 44942 10834 44994
rect 19742 44942 19794 44994
rect 24334 44942 24386 44994
rect 27918 44942 27970 44994
rect 28590 44942 28642 44994
rect 30046 44942 30098 44994
rect 37214 44942 37266 44994
rect 37774 44942 37826 44994
rect 40014 44942 40066 44994
rect 41582 44942 41634 44994
rect 5406 44830 5458 44882
rect 23886 44830 23938 44882
rect 28478 44830 28530 44882
rect 29486 44830 29538 44882
rect 31390 44830 31442 44882
rect 32062 44830 32114 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 30158 44494 30210 44546
rect 40014 44494 40066 44546
rect 40238 44494 40290 44546
rect 1822 44382 1874 44434
rect 28814 44382 28866 44434
rect 30270 44382 30322 44434
rect 31166 44382 31218 44434
rect 31950 44382 32002 44434
rect 33518 44382 33570 44434
rect 10558 44270 10610 44322
rect 11118 44270 11170 44322
rect 12126 44270 12178 44322
rect 15038 44270 15090 44322
rect 15374 44270 15426 44322
rect 31054 44270 31106 44322
rect 19294 44158 19346 44210
rect 32510 44158 32562 44210
rect 58046 44158 58098 44210
rect 7422 44046 7474 44098
rect 8206 44046 8258 44098
rect 11678 44046 11730 44098
rect 14366 44046 14418 44098
rect 17950 44046 18002 44098
rect 18510 44046 18562 44098
rect 18846 44046 18898 44098
rect 31838 44046 31890 44098
rect 32622 44046 32674 44098
rect 33070 44046 33122 44098
rect 40238 44046 40290 44098
rect 57262 44046 57314 44098
rect 57710 44046 57762 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 6190 43710 6242 43762
rect 16158 43710 16210 43762
rect 23438 43710 23490 43762
rect 30606 43710 30658 43762
rect 32510 43710 32562 43762
rect 36766 43710 36818 43762
rect 10222 43598 10274 43650
rect 17726 43598 17778 43650
rect 24334 43598 24386 43650
rect 24894 43598 24946 43650
rect 31614 43598 31666 43650
rect 32062 43598 32114 43650
rect 33966 43598 34018 43650
rect 36878 43598 36930 43650
rect 8542 43486 8594 43538
rect 8878 43486 8930 43538
rect 13022 43486 13074 43538
rect 13582 43486 13634 43538
rect 20302 43486 20354 43538
rect 20974 43486 21026 43538
rect 35086 43486 35138 43538
rect 36654 43486 36706 43538
rect 9662 43374 9714 43426
rect 10782 43374 10834 43426
rect 11342 43374 11394 43426
rect 12126 43374 12178 43426
rect 12686 43374 12738 43426
rect 19854 43374 19906 43426
rect 33854 43374 33906 43426
rect 35534 43374 35586 43426
rect 35982 43374 36034 43426
rect 37102 43374 37154 43426
rect 5406 43262 5458 43314
rect 16718 43262 16770 43314
rect 23998 43262 24050 43314
rect 31502 43262 31554 43314
rect 34750 43262 34802 43314
rect 35086 43262 35138 43314
rect 37326 43262 37378 43314
rect 37550 43262 37602 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 10670 42814 10722 42866
rect 12910 42814 12962 42866
rect 34638 42814 34690 42866
rect 6638 42702 6690 42754
rect 7086 42702 7138 42754
rect 13582 42702 13634 42754
rect 14254 42702 14306 42754
rect 17614 42702 17666 42754
rect 33742 42702 33794 42754
rect 34190 42702 34242 42754
rect 16494 42590 16546 42642
rect 18062 42590 18114 42642
rect 45614 42590 45666 42642
rect 9550 42478 9602 42530
rect 10110 42478 10162 42530
rect 11118 42478 11170 42530
rect 17278 42478 17330 42530
rect 36206 42478 36258 42530
rect 45502 42478 45554 42530
rect 46062 42478 46114 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 2158 42142 2210 42194
rect 23214 42142 23266 42194
rect 10670 42030 10722 42082
rect 1822 41918 1874 41970
rect 15038 41918 15090 41970
rect 20078 41918 20130 41970
rect 20750 41918 20802 41970
rect 24670 41918 24722 41970
rect 15486 41806 15538 41858
rect 19630 41806 19682 41858
rect 24222 41806 24274 41858
rect 23774 41694 23826 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 1822 41246 1874 41298
rect 11006 41246 11058 41298
rect 28814 41246 28866 41298
rect 34190 41246 34242 41298
rect 35534 41246 35586 41298
rect 36430 41246 36482 41298
rect 37886 41246 37938 41298
rect 42814 41246 42866 41298
rect 9774 41134 9826 41186
rect 10334 41134 10386 41186
rect 16718 41134 16770 41186
rect 21534 41134 21586 41186
rect 42142 41134 42194 41186
rect 42590 41134 42642 41186
rect 42926 41134 42978 41186
rect 17390 41022 17442 41074
rect 29598 41022 29650 41074
rect 29822 41022 29874 41074
rect 33630 41022 33682 41074
rect 33742 41022 33794 41074
rect 35982 41022 36034 41074
rect 41806 41022 41858 41074
rect 41918 41022 41970 41074
rect 43262 41022 43314 41074
rect 57262 41022 57314 41074
rect 58046 41022 58098 41074
rect 6638 40910 6690 40962
rect 7422 40910 7474 40962
rect 11342 40910 11394 40962
rect 29710 40910 29762 40962
rect 33406 40910 33458 40962
rect 35086 40910 35138 40962
rect 37550 40910 37602 40962
rect 43822 40910 43874 40962
rect 57710 40910 57762 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 22206 40574 22258 40626
rect 22766 40574 22818 40626
rect 23662 40574 23714 40626
rect 25902 40574 25954 40626
rect 26350 40574 26402 40626
rect 26798 40574 26850 40626
rect 28366 40574 28418 40626
rect 30046 40574 30098 40626
rect 31390 40574 31442 40626
rect 32062 40574 32114 40626
rect 32622 40574 32674 40626
rect 34862 40574 34914 40626
rect 35758 40574 35810 40626
rect 35870 40574 35922 40626
rect 40686 40574 40738 40626
rect 42478 40574 42530 40626
rect 42702 40574 42754 40626
rect 10558 40462 10610 40514
rect 18622 40462 18674 40514
rect 27470 40462 27522 40514
rect 27806 40462 27858 40514
rect 31054 40462 31106 40514
rect 31166 40462 31218 40514
rect 38782 40462 38834 40514
rect 40014 40462 40066 40514
rect 47630 40462 47682 40514
rect 19070 40350 19122 40402
rect 19742 40350 19794 40402
rect 23214 40350 23266 40402
rect 27918 40350 27970 40402
rect 30494 40350 30546 40402
rect 34302 40350 34354 40402
rect 35982 40350 36034 40402
rect 36206 40350 36258 40402
rect 37550 40350 37602 40402
rect 37886 40350 37938 40402
rect 38558 40350 38610 40402
rect 41470 40350 41522 40402
rect 42142 40350 42194 40402
rect 43150 40350 43202 40402
rect 47518 40350 47570 40402
rect 47854 40350 47906 40402
rect 27358 40238 27410 40290
rect 31838 40238 31890 40290
rect 32062 40238 32114 40290
rect 35086 40238 35138 40290
rect 36654 40238 36706 40290
rect 39902 40238 39954 40290
rect 40238 40238 40290 40290
rect 48190 40238 48242 40290
rect 34750 40126 34802 40178
rect 36430 40126 36482 40178
rect 37214 40126 37266 40178
rect 42814 40126 42866 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 20078 39790 20130 39842
rect 33854 39790 33906 39842
rect 40574 39790 40626 39842
rect 20638 39678 20690 39730
rect 27246 39678 27298 39730
rect 28702 39678 28754 39730
rect 37438 39678 37490 39730
rect 38334 39678 38386 39730
rect 41134 39678 41186 39730
rect 42030 39678 42082 39730
rect 42478 39678 42530 39730
rect 16606 39566 16658 39618
rect 17054 39566 17106 39618
rect 21534 39566 21586 39618
rect 28366 39566 28418 39618
rect 28478 39566 28530 39618
rect 31838 39566 31890 39618
rect 35086 39566 35138 39618
rect 35646 39566 35698 39618
rect 38110 39566 38162 39618
rect 38558 39566 38610 39618
rect 39902 39566 39954 39618
rect 40462 39566 40514 39618
rect 47518 39566 47570 39618
rect 48302 39566 48354 39618
rect 28814 39454 28866 39506
rect 31278 39454 31330 39506
rect 31502 39454 31554 39506
rect 32286 39454 32338 39506
rect 33742 39454 33794 39506
rect 34750 39454 34802 39506
rect 34862 39454 34914 39506
rect 36206 39454 36258 39506
rect 38782 39454 38834 39506
rect 39230 39454 39282 39506
rect 40574 39454 40626 39506
rect 47294 39454 47346 39506
rect 48750 39454 48802 39506
rect 48974 39454 49026 39506
rect 19518 39342 19570 39394
rect 26350 39342 26402 39394
rect 26798 39342 26850 39394
rect 27806 39342 27858 39394
rect 31614 39342 31666 39394
rect 33182 39342 33234 39394
rect 35758 39342 35810 39394
rect 35982 39342 36034 39394
rect 36318 39342 36370 39394
rect 36654 39342 36706 39394
rect 41582 39342 41634 39394
rect 46734 39342 46786 39394
rect 47854 39342 47906 39394
rect 48526 39342 48578 39394
rect 49422 39342 49474 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2158 39006 2210 39058
rect 20414 39006 20466 39058
rect 27582 39006 27634 39058
rect 30942 39006 30994 39058
rect 34974 39006 35026 39058
rect 35422 39006 35474 39058
rect 35758 39006 35810 39058
rect 36430 39006 36482 39058
rect 39230 39006 39282 39058
rect 44158 39006 44210 39058
rect 45278 39006 45330 39058
rect 45502 39006 45554 39058
rect 46622 39006 46674 39058
rect 27022 38894 27074 38946
rect 39118 38894 39170 38946
rect 40574 38894 40626 38946
rect 50766 38894 50818 38946
rect 51326 38894 51378 38946
rect 1822 38782 1874 38834
rect 38558 38782 38610 38834
rect 39006 38782 39058 38834
rect 40686 38782 40738 38834
rect 45390 38782 45442 38834
rect 45950 38782 46002 38834
rect 3838 38670 3890 38722
rect 4398 38670 4450 38722
rect 13134 38670 13186 38722
rect 13694 38670 13746 38722
rect 14702 38670 14754 38722
rect 15150 38670 15202 38722
rect 34414 38670 34466 38722
rect 41582 38670 41634 38722
rect 41918 38670 41970 38722
rect 44606 38670 44658 38722
rect 45726 38670 45778 38722
rect 3950 38558 4002 38610
rect 26910 38558 26962 38610
rect 46174 38558 46226 38610
rect 50878 38558 50930 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 26574 38222 26626 38274
rect 1822 38110 1874 38162
rect 12014 38110 12066 38162
rect 24558 38110 24610 38162
rect 34414 38110 34466 38162
rect 35086 38110 35138 38162
rect 41134 38110 41186 38162
rect 41694 38110 41746 38162
rect 14254 37998 14306 38050
rect 14590 37998 14642 38050
rect 25566 37998 25618 38050
rect 26126 37998 26178 38050
rect 30830 37998 30882 38050
rect 31166 37998 31218 38050
rect 31502 37998 31554 38050
rect 32846 37998 32898 38050
rect 33518 37998 33570 38050
rect 33966 37998 34018 38050
rect 35310 37998 35362 38050
rect 39454 37998 39506 38050
rect 39790 37998 39842 38050
rect 40910 37998 40962 38050
rect 42142 37998 42194 38050
rect 12910 37886 12962 37938
rect 14030 37886 14082 37938
rect 15150 37886 15202 37938
rect 25678 37886 25730 37938
rect 25902 37886 25954 37938
rect 30158 37886 30210 37938
rect 30382 37886 30434 37938
rect 35982 37886 36034 37938
rect 36654 37886 36706 37938
rect 39118 37886 39170 37938
rect 40238 37886 40290 37938
rect 58046 37886 58098 37938
rect 12686 37774 12738 37826
rect 12798 37774 12850 37826
rect 13918 37774 13970 37826
rect 15038 37774 15090 37826
rect 15598 37774 15650 37826
rect 18510 37774 18562 37826
rect 19070 37774 19122 37826
rect 24110 37774 24162 37826
rect 25006 37774 25058 37826
rect 26910 37774 26962 37826
rect 27358 37774 27410 37826
rect 30606 37774 30658 37826
rect 31390 37774 31442 37826
rect 31950 37774 32002 37826
rect 32398 37774 32450 37826
rect 32958 37774 33010 37826
rect 33182 37774 33234 37826
rect 36542 37774 36594 37826
rect 39454 37774 39506 37826
rect 57262 37774 57314 37826
rect 57710 37774 57762 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 10894 37438 10946 37490
rect 13358 37438 13410 37490
rect 16942 37438 16994 37490
rect 19854 37438 19906 37490
rect 20526 37438 20578 37490
rect 27358 37438 27410 37490
rect 32622 37438 32674 37490
rect 36206 37438 36258 37490
rect 12014 37326 12066 37378
rect 17726 37326 17778 37378
rect 25006 37326 25058 37378
rect 25790 37326 25842 37378
rect 27246 37326 27298 37378
rect 30942 37326 30994 37378
rect 31502 37326 31554 37378
rect 40462 37326 40514 37378
rect 40686 37326 40738 37378
rect 12574 37214 12626 37266
rect 12798 37214 12850 37266
rect 13246 37214 13298 37266
rect 13470 37214 13522 37266
rect 19294 37214 19346 37266
rect 19742 37214 19794 37266
rect 19966 37214 20018 37266
rect 20974 37214 21026 37266
rect 25678 37214 25730 37266
rect 28814 37214 28866 37266
rect 29150 37214 29202 37266
rect 41470 37214 41522 37266
rect 49646 37214 49698 37266
rect 49982 37214 50034 37266
rect 5070 37102 5122 37154
rect 8766 37102 8818 37154
rect 11454 37102 11506 37154
rect 13022 37102 13074 37154
rect 14030 37102 14082 37154
rect 14478 37102 14530 37154
rect 14926 37102 14978 37154
rect 15374 37102 15426 37154
rect 16494 37102 16546 37154
rect 18510 37102 18562 37154
rect 19518 37102 19570 37154
rect 26574 37102 26626 37154
rect 39790 37102 39842 37154
rect 40574 37102 40626 37154
rect 49534 37102 49586 37154
rect 50990 37102 51042 37154
rect 11902 36990 11954 37042
rect 17838 36990 17890 37042
rect 19070 36990 19122 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 3838 36654 3890 36706
rect 31054 36654 31106 36706
rect 34078 36654 34130 36706
rect 41358 36654 41410 36706
rect 42478 36654 42530 36706
rect 49534 36654 49586 36706
rect 4062 36542 4114 36594
rect 4510 36542 4562 36594
rect 5630 36542 5682 36594
rect 8094 36542 8146 36594
rect 8878 36542 8930 36594
rect 11454 36542 11506 36594
rect 12686 36542 12738 36594
rect 13694 36542 13746 36594
rect 14590 36542 14642 36594
rect 16942 36542 16994 36594
rect 17390 36542 17442 36594
rect 19070 36542 19122 36594
rect 19854 36542 19906 36594
rect 20414 36542 20466 36594
rect 24894 36542 24946 36594
rect 27134 36542 27186 36594
rect 30494 36542 30546 36594
rect 32286 36542 32338 36594
rect 32734 36542 32786 36594
rect 34414 36542 34466 36594
rect 34862 36542 34914 36594
rect 40798 36542 40850 36594
rect 41582 36542 41634 36594
rect 42142 36542 42194 36594
rect 42926 36542 42978 36594
rect 43486 36542 43538 36594
rect 4398 36430 4450 36482
rect 6414 36430 6466 36482
rect 7310 36430 7362 36482
rect 7534 36430 7586 36482
rect 7870 36430 7922 36482
rect 8206 36430 8258 36482
rect 11902 36430 11954 36482
rect 12126 36430 12178 36482
rect 12462 36430 12514 36482
rect 14142 36430 14194 36482
rect 19182 36430 19234 36482
rect 19406 36430 19458 36482
rect 19630 36430 19682 36482
rect 25230 36430 25282 36482
rect 25454 36430 25506 36482
rect 25678 36430 25730 36482
rect 30606 36430 30658 36482
rect 30718 36430 30770 36482
rect 31278 36430 31330 36482
rect 32174 36430 32226 36482
rect 33518 36430 33570 36482
rect 34078 36430 34130 36482
rect 41134 36430 41186 36482
rect 1822 36318 1874 36370
rect 8990 36318 9042 36370
rect 9214 36318 9266 36370
rect 12798 36318 12850 36370
rect 15934 36318 15986 36370
rect 16158 36318 16210 36370
rect 18286 36318 18338 36370
rect 23550 36318 23602 36370
rect 24110 36318 24162 36370
rect 40014 36318 40066 36370
rect 42254 36318 42306 36370
rect 2158 36206 2210 36258
rect 4510 36206 4562 36258
rect 4734 36206 4786 36258
rect 6862 36206 6914 36258
rect 7982 36206 8034 36258
rect 9774 36206 9826 36258
rect 10110 36206 10162 36258
rect 10558 36206 10610 36258
rect 12574 36206 12626 36258
rect 15374 36206 15426 36258
rect 16046 36206 16098 36258
rect 16830 36206 16882 36258
rect 17838 36206 17890 36258
rect 18958 36206 19010 36258
rect 22878 36206 22930 36258
rect 23438 36206 23490 36258
rect 24782 36206 24834 36258
rect 25006 36206 25058 36258
rect 26238 36206 26290 36258
rect 26574 36206 26626 36258
rect 29710 36206 29762 36258
rect 30382 36206 30434 36258
rect 39566 36206 39618 36258
rect 40686 36206 40738 36258
rect 40910 36206 40962 36258
rect 49310 36206 49362 36258
rect 49422 36206 49474 36258
rect 49982 36206 50034 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 5294 35870 5346 35922
rect 8206 35870 8258 35922
rect 14142 35870 14194 35922
rect 14702 35870 14754 35922
rect 16158 35870 16210 35922
rect 17166 35870 17218 35922
rect 17838 35870 17890 35922
rect 1710 35758 1762 35810
rect 8766 35758 8818 35810
rect 8878 35758 8930 35810
rect 9774 35758 9826 35810
rect 12910 35758 12962 35810
rect 14254 35758 14306 35810
rect 15374 35758 15426 35810
rect 9102 35646 9154 35698
rect 10110 35646 10162 35698
rect 16046 35646 16098 35698
rect 16270 35646 16322 35698
rect 16494 35646 16546 35698
rect 16718 35646 16770 35698
rect 16942 35646 16994 35698
rect 10446 35534 10498 35586
rect 11342 35534 11394 35586
rect 11790 35534 11842 35586
rect 13358 35534 13410 35586
rect 18734 35870 18786 35922
rect 20078 35870 20130 35922
rect 32846 35870 32898 35922
rect 35982 35870 36034 35922
rect 39678 35870 39730 35922
rect 44718 35870 44770 35922
rect 45166 35870 45218 35922
rect 45950 35870 46002 35922
rect 46062 35870 46114 35922
rect 18286 35758 18338 35810
rect 29710 35758 29762 35810
rect 33630 35758 33682 35810
rect 35086 35758 35138 35810
rect 35646 35758 35698 35810
rect 35758 35758 35810 35810
rect 38222 35758 38274 35810
rect 39566 35758 39618 35810
rect 45838 35758 45890 35810
rect 47294 35758 47346 35810
rect 49534 35758 49586 35810
rect 19294 35646 19346 35698
rect 19854 35646 19906 35698
rect 19966 35646 20018 35698
rect 20190 35646 20242 35698
rect 32398 35646 32450 35698
rect 33742 35646 33794 35698
rect 34414 35646 34466 35698
rect 34974 35646 35026 35698
rect 39790 35646 39842 35698
rect 46286 35646 46338 35698
rect 46510 35646 46562 35698
rect 50094 35646 50146 35698
rect 50878 35646 50930 35698
rect 51886 35646 51938 35698
rect 31502 35534 31554 35586
rect 36318 35534 36370 35586
rect 38670 35534 38722 35586
rect 40014 35534 40066 35586
rect 41806 35534 41858 35586
rect 51326 35534 51378 35586
rect 17166 35422 17218 35474
rect 19518 35422 19570 35474
rect 40238 35422 40290 35474
rect 40462 35422 40514 35474
rect 46734 35422 46786 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19406 35086 19458 35138
rect 23662 35086 23714 35138
rect 24558 35086 24610 35138
rect 24782 35086 24834 35138
rect 29598 35086 29650 35138
rect 8990 34974 9042 35026
rect 12238 34974 12290 35026
rect 15150 34974 15202 35026
rect 15934 34974 15986 35026
rect 16942 34974 16994 35026
rect 21870 34974 21922 35026
rect 22430 34974 22482 35026
rect 22990 34974 23042 35026
rect 25454 34974 25506 35026
rect 26686 34974 26738 35026
rect 33294 34974 33346 35026
rect 35646 34974 35698 35026
rect 44718 34974 44770 35026
rect 46062 34974 46114 35026
rect 56254 34974 56306 35026
rect 57822 34974 57874 35026
rect 11678 34862 11730 34914
rect 15486 34862 15538 34914
rect 17614 34862 17666 34914
rect 17950 34862 18002 34914
rect 22094 34862 22146 34914
rect 25006 34862 25058 34914
rect 25230 34862 25282 34914
rect 26350 34862 26402 34914
rect 34526 34862 34578 34914
rect 34862 34862 34914 34914
rect 35086 34862 35138 34914
rect 40238 34862 40290 34914
rect 40462 34862 40514 34914
rect 45838 34862 45890 34914
rect 56814 34862 56866 34914
rect 9550 34750 9602 34802
rect 10222 34750 10274 34802
rect 10558 34750 10610 34802
rect 10782 34750 10834 34802
rect 18510 34750 18562 34802
rect 19070 34750 19122 34802
rect 25454 34750 25506 34802
rect 29710 34750 29762 34802
rect 46174 34750 46226 34802
rect 9662 34638 9714 34690
rect 10334 34638 10386 34690
rect 19294 34638 19346 34690
rect 19854 34638 19906 34690
rect 20414 34638 20466 34690
rect 20862 34638 20914 34690
rect 21758 34638 21810 34690
rect 21982 34638 22034 34690
rect 23326 34638 23378 34690
rect 23774 34638 23826 34690
rect 24222 34638 24274 34690
rect 25678 34638 25730 34690
rect 30158 34638 30210 34690
rect 34862 34638 34914 34690
rect 36094 34638 36146 34690
rect 39118 34638 39170 34690
rect 39902 34638 39954 34690
rect 46622 34638 46674 34690
rect 50318 34638 50370 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 8542 34302 8594 34354
rect 10558 34302 10610 34354
rect 34414 34302 34466 34354
rect 34526 34302 34578 34354
rect 36094 34302 36146 34354
rect 36542 34302 36594 34354
rect 37438 34302 37490 34354
rect 45166 34302 45218 34354
rect 45838 34302 45890 34354
rect 45950 34302 46002 34354
rect 4734 34190 4786 34242
rect 7982 34190 8034 34242
rect 8094 34190 8146 34242
rect 10446 34190 10498 34242
rect 36766 34190 36818 34242
rect 5070 34078 5122 34130
rect 9998 34078 10050 34130
rect 10670 34078 10722 34130
rect 11230 34078 11282 34130
rect 34638 34078 34690 34130
rect 35086 34078 35138 34130
rect 4958 33966 5010 34018
rect 5518 33966 5570 34018
rect 9774 33966 9826 34018
rect 10222 33966 10274 34018
rect 11678 33966 11730 34018
rect 19854 33966 19906 34018
rect 20414 33966 20466 34018
rect 26574 33966 26626 34018
rect 27022 33966 27074 34018
rect 33854 33966 33906 34018
rect 35646 33966 35698 34018
rect 19966 33854 20018 33906
rect 36206 33854 36258 33906
rect 36990 33966 37042 34018
rect 37886 33966 37938 34018
rect 46622 33966 46674 34018
rect 37438 33854 37490 33906
rect 37998 33854 38050 33906
rect 46062 33854 46114 33906
rect 46286 33854 46338 33906
rect 46622 33854 46674 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 26462 33518 26514 33570
rect 32622 33518 32674 33570
rect 34750 33518 34802 33570
rect 34974 33518 35026 33570
rect 35198 33518 35250 33570
rect 38334 33518 38386 33570
rect 11454 33406 11506 33458
rect 11902 33406 11954 33458
rect 17278 33406 17330 33458
rect 23998 33406 24050 33458
rect 24446 33406 24498 33458
rect 25454 33406 25506 33458
rect 30270 33406 30322 33458
rect 36318 33406 36370 33458
rect 40014 33406 40066 33458
rect 42030 33406 42082 33458
rect 42478 33406 42530 33458
rect 49534 33406 49586 33458
rect 16158 33294 16210 33346
rect 16718 33294 16770 33346
rect 25790 33294 25842 33346
rect 26126 33294 26178 33346
rect 35422 33294 35474 33346
rect 36094 33294 36146 33346
rect 36766 33294 36818 33346
rect 37998 33294 38050 33346
rect 38558 33294 38610 33346
rect 41918 33294 41970 33346
rect 25566 33182 25618 33234
rect 26798 33182 26850 33234
rect 27022 33182 27074 33234
rect 27134 33182 27186 33234
rect 27806 33182 27858 33234
rect 28254 33182 28306 33234
rect 29598 33182 29650 33234
rect 29710 33182 29762 33234
rect 32286 33182 32338 33234
rect 36542 33182 36594 33234
rect 25006 33070 25058 33122
rect 27694 33070 27746 33122
rect 28926 33070 28978 33122
rect 29934 33070 29986 33122
rect 31726 33070 31778 33122
rect 32510 33070 32562 33122
rect 33070 33070 33122 33122
rect 34302 33070 34354 33122
rect 37662 33070 37714 33122
rect 37774 33070 37826 33122
rect 37886 33070 37938 33122
rect 39006 33070 39058 33122
rect 39566 33070 39618 33122
rect 50094 33070 50146 33122
rect 50542 33070 50594 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 3502 32734 3554 32786
rect 9998 32734 10050 32786
rect 11454 32734 11506 32786
rect 12238 32734 12290 32786
rect 21646 32734 21698 32786
rect 22542 32734 22594 32786
rect 26350 32734 26402 32786
rect 27246 32734 27298 32786
rect 27358 32734 27410 32786
rect 27470 32734 27522 32786
rect 28590 32734 28642 32786
rect 33966 32734 34018 32786
rect 34526 32734 34578 32786
rect 34750 32734 34802 32786
rect 35534 32734 35586 32786
rect 37214 32734 37266 32786
rect 38222 32734 38274 32786
rect 38894 32734 38946 32786
rect 39566 32734 39618 32786
rect 11566 32622 11618 32674
rect 12462 32622 12514 32674
rect 35310 32622 35362 32674
rect 37326 32622 37378 32674
rect 42702 32622 42754 32674
rect 3054 32510 3106 32562
rect 9886 32510 9938 32562
rect 10110 32510 10162 32562
rect 10334 32510 10386 32562
rect 10782 32510 10834 32562
rect 11230 32510 11282 32562
rect 12014 32510 12066 32562
rect 12574 32510 12626 32562
rect 21422 32510 21474 32562
rect 21758 32510 21810 32562
rect 22206 32510 22258 32562
rect 22654 32510 22706 32562
rect 22878 32510 22930 32562
rect 26014 32510 26066 32562
rect 26238 32510 26290 32562
rect 26686 32510 26738 32562
rect 27582 32510 27634 32562
rect 34414 32510 34466 32562
rect 35198 32510 35250 32562
rect 42142 32510 42194 32562
rect 2046 32398 2098 32450
rect 13134 32398 13186 32450
rect 23326 32398 23378 32450
rect 23774 32398 23826 32450
rect 24894 32398 24946 32450
rect 35870 32398 35922 32450
rect 36318 32398 36370 32450
rect 38110 32398 38162 32450
rect 40126 32398 40178 32450
rect 40686 32398 40738 32450
rect 10558 32286 10610 32338
rect 27918 32286 27970 32338
rect 28142 32286 28194 32338
rect 38446 32286 38498 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 11006 31838 11058 31890
rect 16046 31838 16098 31890
rect 17166 31838 17218 31890
rect 17502 31838 17554 31890
rect 23662 31838 23714 31890
rect 26910 31838 26962 31890
rect 27246 31838 27298 31890
rect 30494 31838 30546 31890
rect 35758 31838 35810 31890
rect 39230 31838 39282 31890
rect 39902 31838 39954 31890
rect 36878 31726 36930 31778
rect 38110 31726 38162 31778
rect 38558 31726 38610 31778
rect 39118 31726 39170 31778
rect 41806 31726 41858 31778
rect 11902 31614 11954 31666
rect 16606 31614 16658 31666
rect 17054 31614 17106 31666
rect 23886 31614 23938 31666
rect 30830 31614 30882 31666
rect 37886 31614 37938 31666
rect 37998 31614 38050 31666
rect 39454 31614 39506 31666
rect 41246 31614 41298 31666
rect 11678 31502 11730 31554
rect 11790 31502 11842 31554
rect 12350 31502 12402 31554
rect 16830 31502 16882 31554
rect 18062 31502 18114 31554
rect 21982 31502 22034 31554
rect 23662 31502 23714 31554
rect 24334 31502 24386 31554
rect 24782 31502 24834 31554
rect 30606 31502 30658 31554
rect 31278 31502 31330 31554
rect 31726 31502 31778 31554
rect 34078 31502 34130 31554
rect 40350 31502 40402 31554
rect 41358 31502 41410 31554
rect 58046 31502 58098 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 10446 31166 10498 31218
rect 10894 31166 10946 31218
rect 29486 31166 29538 31218
rect 39902 31166 39954 31218
rect 40014 31166 40066 31218
rect 40574 31166 40626 31218
rect 12014 31054 12066 31106
rect 12126 31054 12178 31106
rect 12686 31054 12738 31106
rect 5518 30942 5570 30994
rect 11342 30942 11394 30994
rect 13134 30942 13186 30994
rect 28926 30942 28978 30994
rect 4734 30830 4786 30882
rect 5182 30830 5234 30882
rect 5966 30830 6018 30882
rect 13022 30830 13074 30882
rect 19070 30830 19122 30882
rect 28142 30830 28194 30882
rect 28702 30830 28754 30882
rect 37438 30830 37490 30882
rect 40126 30830 40178 30882
rect 41582 30830 41634 30882
rect 5518 30718 5570 30770
rect 12014 30718 12066 30770
rect 28590 30718 28642 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 8654 30382 8706 30434
rect 9214 30382 9266 30434
rect 9438 30382 9490 30434
rect 19182 30382 19234 30434
rect 32062 30382 32114 30434
rect 5742 30270 5794 30322
rect 6078 30270 6130 30322
rect 17726 30270 17778 30322
rect 6526 30158 6578 30210
rect 9662 30158 9714 30210
rect 9886 30158 9938 30210
rect 9998 30158 10050 30210
rect 10670 30158 10722 30210
rect 12350 30158 12402 30210
rect 12798 30158 12850 30210
rect 13582 30158 13634 30210
rect 13918 30158 13970 30210
rect 14366 30158 14418 30210
rect 16046 30158 16098 30210
rect 17166 30158 17218 30210
rect 17950 30158 18002 30210
rect 18286 30158 18338 30210
rect 18622 30158 18674 30210
rect 19630 30158 19682 30210
rect 19854 30158 19906 30210
rect 20190 30158 20242 30210
rect 21646 30158 21698 30210
rect 1822 30046 1874 30098
rect 2158 30046 2210 30098
rect 5966 30046 6018 30098
rect 8318 30046 8370 30098
rect 8542 30046 8594 30098
rect 10110 30046 10162 30098
rect 12238 30046 12290 30098
rect 13806 30046 13858 30098
rect 14926 30046 14978 30098
rect 15486 30046 15538 30098
rect 19966 30046 20018 30098
rect 20862 30046 20914 30098
rect 32622 30046 32674 30098
rect 7758 29934 7810 29986
rect 11342 29934 11394 29986
rect 16830 29934 16882 29986
rect 18398 29934 18450 29986
rect 18510 29934 18562 29986
rect 31166 29934 31218 29986
rect 31614 29934 31666 29986
rect 32174 29934 32226 29986
rect 32398 29934 32450 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 1822 29598 1874 29650
rect 8990 29598 9042 29650
rect 10894 29598 10946 29650
rect 11678 29598 11730 29650
rect 14142 29598 14194 29650
rect 17054 29598 17106 29650
rect 17614 29598 17666 29650
rect 19182 29598 19234 29650
rect 20414 29598 20466 29650
rect 24894 29598 24946 29650
rect 25678 29598 25730 29650
rect 34414 29598 34466 29650
rect 57710 29598 57762 29650
rect 12238 29486 12290 29538
rect 18286 29486 18338 29538
rect 19518 29486 19570 29538
rect 26238 29486 26290 29538
rect 10558 29374 10610 29426
rect 10782 29374 10834 29426
rect 11230 29374 11282 29426
rect 18510 29374 18562 29426
rect 18958 29374 19010 29426
rect 22654 29374 22706 29426
rect 23102 29374 23154 29426
rect 23326 29374 23378 29426
rect 33630 29374 33682 29426
rect 58046 29374 58098 29426
rect 18174 29262 18226 29314
rect 22206 29262 22258 29314
rect 23214 29262 23266 29314
rect 23774 29262 23826 29314
rect 24222 29262 24274 29314
rect 32174 29262 32226 29314
rect 32734 29262 32786 29314
rect 33742 29262 33794 29314
rect 32846 29150 32898 29202
rect 33966 29150 34018 29202
rect 34190 29150 34242 29202
rect 34414 29150 34466 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 11342 28814 11394 28866
rect 11566 28814 11618 28866
rect 12014 28814 12066 28866
rect 12350 28814 12402 28866
rect 16606 28814 16658 28866
rect 34190 28814 34242 28866
rect 34526 28814 34578 28866
rect 11342 28702 11394 28754
rect 12574 28702 12626 28754
rect 13582 28702 13634 28754
rect 15822 28702 15874 28754
rect 16382 28702 16434 28754
rect 16942 28702 16994 28754
rect 17726 28702 17778 28754
rect 19406 28702 19458 28754
rect 23550 28702 23602 28754
rect 26462 28702 26514 28754
rect 27918 28702 27970 28754
rect 28478 28702 28530 28754
rect 33294 28702 33346 28754
rect 34190 28702 34242 28754
rect 34638 28702 34690 28754
rect 35758 28702 35810 28754
rect 58158 28702 58210 28754
rect 18174 28590 18226 28642
rect 18286 28590 18338 28642
rect 18734 28590 18786 28642
rect 18958 28590 19010 28642
rect 23102 28590 23154 28642
rect 23438 28590 23490 28642
rect 24222 28590 24274 28642
rect 24670 28590 24722 28642
rect 27470 28590 27522 28642
rect 35982 28590 36034 28642
rect 38110 28590 38162 28642
rect 38558 28590 38610 28642
rect 39566 28590 39618 28642
rect 39902 28590 39954 28642
rect 40462 28590 40514 28642
rect 42254 28590 42306 28642
rect 18510 28478 18562 28530
rect 27022 28478 27074 28530
rect 35310 28478 35362 28530
rect 35534 28478 35586 28530
rect 39118 28478 39170 28530
rect 39342 28478 39394 28530
rect 41358 28478 41410 28530
rect 22990 28366 23042 28418
rect 35422 28366 35474 28418
rect 39902 28366 39954 28418
rect 41694 28366 41746 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 6078 28030 6130 28082
rect 7310 28030 7362 28082
rect 10894 28030 10946 28082
rect 12014 28030 12066 28082
rect 12910 28030 12962 28082
rect 17726 28030 17778 28082
rect 23326 28030 23378 28082
rect 28702 28030 28754 28082
rect 29262 28030 29314 28082
rect 23214 27918 23266 27970
rect 23774 27918 23826 27970
rect 24222 27918 24274 27970
rect 28814 27918 28866 27970
rect 6302 27806 6354 27858
rect 6750 27806 6802 27858
rect 10558 27806 10610 27858
rect 10782 27806 10834 27858
rect 11006 27806 11058 27858
rect 11566 27806 11618 27858
rect 23550 27806 23602 27858
rect 6078 27694 6130 27746
rect 10110 27694 10162 27746
rect 24670 27694 24722 27746
rect 10334 27582 10386 27634
rect 28702 27582 28754 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 18734 27246 18786 27298
rect 25342 27246 25394 27298
rect 34078 27246 34130 27298
rect 3502 27134 3554 27186
rect 11454 27134 11506 27186
rect 17838 27134 17890 27186
rect 18286 27134 18338 27186
rect 20190 27134 20242 27186
rect 24558 27134 24610 27186
rect 26014 27134 26066 27186
rect 29486 27134 29538 27186
rect 31278 27134 31330 27186
rect 3054 27022 3106 27074
rect 11678 27022 11730 27074
rect 12126 27022 12178 27074
rect 17390 27022 17442 27074
rect 19182 27022 19234 27074
rect 19406 27022 19458 27074
rect 19630 27022 19682 27074
rect 22878 27022 22930 27074
rect 23326 27022 23378 27074
rect 23550 27022 23602 27074
rect 24446 27022 24498 27074
rect 24782 27022 24834 27074
rect 25118 27022 25170 27074
rect 27694 27022 27746 27074
rect 28030 27022 28082 27074
rect 31726 27022 31778 27074
rect 32734 27022 32786 27074
rect 33294 27022 33346 27074
rect 33742 27022 33794 27074
rect 2158 26910 2210 26962
rect 11342 26910 11394 26962
rect 19518 26910 19570 26962
rect 24670 26910 24722 26962
rect 26462 26910 26514 26962
rect 27022 26910 27074 26962
rect 28590 26910 28642 26962
rect 32622 26910 32674 26962
rect 23214 26798 23266 26850
rect 28478 26798 28530 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 10222 26462 10274 26514
rect 11342 26462 11394 26514
rect 12462 26462 12514 26514
rect 23662 26462 23714 26514
rect 23998 26462 24050 26514
rect 24558 26462 24610 26514
rect 25678 26462 25730 26514
rect 27246 26462 27298 26514
rect 27806 26462 27858 26514
rect 32174 26462 32226 26514
rect 42030 26462 42082 26514
rect 42702 26462 42754 26514
rect 12014 26350 12066 26402
rect 27022 26350 27074 26402
rect 41582 26350 41634 26402
rect 10782 26238 10834 26290
rect 41918 26238 41970 26290
rect 42142 26238 42194 26290
rect 27358 26126 27410 26178
rect 43038 26126 43090 26178
rect 11902 26014 11954 26066
rect 42366 26014 42418 26066
rect 43038 26014 43090 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 22542 25678 22594 25730
rect 24110 25678 24162 25730
rect 9774 25566 9826 25618
rect 10670 25566 10722 25618
rect 11566 25566 11618 25618
rect 22430 25566 22482 25618
rect 22990 25566 23042 25618
rect 56254 25566 56306 25618
rect 57822 25566 57874 25618
rect 10894 25454 10946 25506
rect 56814 25454 56866 25506
rect 9774 25342 9826 25394
rect 9998 25342 10050 25394
rect 23998 25342 24050 25394
rect 24110 25230 24162 25282
rect 24670 25230 24722 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 9774 24894 9826 24946
rect 10334 24894 10386 24946
rect 10782 24894 10834 24946
rect 19742 24894 19794 24946
rect 21758 24894 21810 24946
rect 22318 24894 22370 24946
rect 23214 24894 23266 24946
rect 24670 24894 24722 24946
rect 24782 24894 24834 24946
rect 26910 24894 26962 24946
rect 27470 24894 27522 24946
rect 27806 24894 27858 24946
rect 28254 24894 28306 24946
rect 28366 24894 28418 24946
rect 28590 24894 28642 24946
rect 10894 24782 10946 24834
rect 11342 24782 11394 24834
rect 12238 24782 12290 24834
rect 28814 24782 28866 24834
rect 11118 24670 11170 24722
rect 24222 24670 24274 24722
rect 24446 24670 24498 24722
rect 11790 24558 11842 24610
rect 19630 24558 19682 24610
rect 22430 24558 22482 24610
rect 23662 24558 23714 24610
rect 9774 24446 9826 24498
rect 10670 24446 10722 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3614 23998 3666 24050
rect 18174 23998 18226 24050
rect 18622 23998 18674 24050
rect 25118 23998 25170 24050
rect 26350 23998 26402 24050
rect 3054 23886 3106 23938
rect 17166 23886 17218 23938
rect 17390 23886 17442 23938
rect 22766 23886 22818 23938
rect 24334 23886 24386 23938
rect 2158 23774 2210 23826
rect 17726 23774 17778 23826
rect 23214 23774 23266 23826
rect 24222 23774 24274 23826
rect 21646 23662 21698 23714
rect 22094 23662 22146 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 11342 23326 11394 23378
rect 18062 23326 18114 23378
rect 18846 23326 18898 23378
rect 19182 23326 19234 23378
rect 21198 23326 21250 23378
rect 22094 23326 22146 23378
rect 23550 23326 23602 23378
rect 9774 23214 9826 23266
rect 17950 23214 18002 23266
rect 22990 23214 23042 23266
rect 57710 23214 57762 23266
rect 10446 23102 10498 23154
rect 17838 23102 17890 23154
rect 18398 23102 18450 23154
rect 22318 23102 22370 23154
rect 22766 23102 22818 23154
rect 23102 23102 23154 23154
rect 58046 23102 58098 23154
rect 10670 22990 10722 23042
rect 11678 22990 11730 23042
rect 16942 22990 16994 23042
rect 21646 22990 21698 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 11006 22542 11058 22594
rect 9438 22430 9490 22482
rect 11790 22430 11842 22482
rect 58158 22430 58210 22482
rect 10110 22318 10162 22370
rect 10334 22318 10386 22370
rect 10558 22318 10610 22370
rect 12238 22318 12290 22370
rect 9998 22206 10050 22258
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 3502 21758 3554 21810
rect 11342 21758 11394 21810
rect 3054 21534 3106 21586
rect 2046 21422 2098 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4286 20862 4338 20914
rect 57710 20638 57762 20690
rect 58046 20638 58098 20690
rect 3726 20526 3778 20578
rect 57262 20526 57314 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 1822 17502 1874 17554
rect 2158 17502 2210 17554
rect 57710 17502 57762 17554
rect 58046 17502 58098 17554
rect 57262 17390 57314 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 1822 17054 1874 17106
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2158 15486 2210 15538
rect 1822 15262 1874 15314
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14590 1874 14642
rect 56366 14590 56418 14642
rect 56814 14478 56866 14530
rect 57710 14366 57762 14418
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 3502 12350 3554 12402
rect 3054 12126 3106 12178
rect 2046 12014 2098 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 56814 11342 56866 11394
rect 57710 11230 57762 11282
rect 56366 11118 56418 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 2158 9214 2210 9266
rect 1822 8990 1874 9042
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 1822 8318 1874 8370
rect 57710 8094 57762 8146
rect 58046 8094 58098 8146
rect 57262 7982 57314 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 3502 6078 3554 6130
rect 58046 5966 58098 6018
rect 3054 5854 3106 5906
rect 2046 5742 2098 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 3614 5182 3666 5234
rect 3054 5070 3106 5122
rect 2158 4958 2210 5010
rect 57262 4958 57314 5010
rect 57710 4958 57762 5010
rect 58046 4958 58098 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 3502 4510 3554 4562
rect 4398 4510 4450 4562
rect 11118 4510 11170 4562
rect 16494 4510 16546 4562
rect 34750 4510 34802 4562
rect 57710 4510 57762 4562
rect 3054 4286 3106 4338
rect 58046 4286 58098 4338
rect 2046 4174 2098 4226
rect 56814 4174 56866 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 15262 3614 15314 3666
rect 16830 3614 16882 3666
rect 18398 3614 18450 3666
rect 32510 3614 32562 3666
rect 35758 3614 35810 3666
rect 44270 3614 44322 3666
rect 45166 3614 45218 3666
rect 4174 3502 4226 3554
rect 10894 3502 10946 3554
rect 16270 3502 16322 3554
rect 17726 3502 17778 3554
rect 33182 3502 33234 3554
rect 35086 3502 35138 3554
rect 45950 3502 46002 3554
rect 56030 3502 56082 3554
rect 56702 3502 56754 3554
rect 3278 3390 3330 3442
rect 5070 3390 5122 3442
rect 5742 3390 5794 3442
rect 9998 3390 10050 3442
rect 20750 3390 20802 3442
rect 21422 3390 21474 3442
rect 23326 3390 23378 3442
rect 23774 3390 23826 3442
rect 29374 3390 29426 3442
rect 29822 3390 29874 3442
rect 34078 3390 34130 3442
rect 41470 3390 41522 3442
rect 41918 3390 41970 3442
rect 48190 3390 48242 3442
rect 49198 3390 49250 3442
rect 50206 3390 50258 3442
rect 50990 3390 51042 3442
rect 57598 3390 57650 3442
rect 6078 3278 6130 3330
rect 11678 3278 11730 3330
rect 21758 3278 21810 3330
rect 24110 3278 24162 3330
rect 27134 3278 27186 3330
rect 30158 3278 30210 3330
rect 42254 3278 42306 3330
rect 48862 3278 48914 3330
rect 50654 3278 50706 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 1960 59304 2184 59800
rect 1960 59220 2212 59304
rect 2268 59276 2660 59332
rect 2268 59220 2324 59276
rect 1960 59200 2324 59220
rect 2156 59164 2324 59200
rect 1820 56420 1876 56430
rect 1820 55186 1876 56364
rect 2604 56194 2660 59276
rect 4648 59304 4872 59800
rect 8008 59304 8232 59800
rect 10696 59304 10920 59800
rect 4648 59200 4900 59304
rect 8008 59200 8260 59304
rect 10696 59220 10948 59304
rect 11004 59276 11396 59332
rect 14056 59304 14280 59800
rect 11004 59220 11060 59276
rect 10696 59200 11060 59220
rect 2604 56142 2606 56194
rect 2658 56142 2660 56194
rect 2604 56130 2660 56142
rect 4844 56196 4900 59200
rect 8204 56308 8260 59200
rect 10892 59164 11060 59200
rect 8316 56308 8372 56318
rect 8204 56306 8372 56308
rect 8204 56254 8318 56306
rect 8370 56254 8372 56306
rect 8204 56252 8372 56254
rect 8316 56242 8372 56252
rect 4844 56130 4900 56140
rect 6076 56196 6132 56206
rect 6076 56102 6132 56140
rect 11340 56194 11396 59276
rect 11340 56142 11342 56194
rect 11394 56142 11396 56194
rect 11340 56130 11396 56142
rect 14028 59200 14280 59304
rect 16744 59304 16968 59800
rect 16744 59220 16996 59304
rect 17052 59276 17780 59332
rect 19432 59304 19656 59800
rect 17052 59220 17108 59276
rect 16744 59200 17108 59220
rect 3500 56082 3556 56094
rect 3500 56030 3502 56082
rect 3554 56030 3556 56082
rect 3500 55972 3556 56030
rect 6972 56084 7028 56094
rect 7532 56084 7588 56094
rect 6972 56082 7588 56084
rect 6972 56030 6974 56082
rect 7026 56030 7534 56082
rect 7586 56030 7588 56082
rect 6972 56028 7588 56030
rect 6972 56018 7028 56028
rect 3500 55906 3556 55916
rect 4060 55972 4116 55982
rect 4060 55878 4116 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 1820 55134 1822 55186
rect 1874 55134 1876 55186
rect 1820 54738 1876 55134
rect 2156 55076 2212 55086
rect 2156 55074 2324 55076
rect 2156 55022 2158 55074
rect 2210 55022 2324 55074
rect 2156 55020 2324 55022
rect 2156 55010 2212 55020
rect 1820 54686 1822 54738
rect 1874 54686 1876 54738
rect 1820 54674 1876 54686
rect 2044 53844 2100 53854
rect 1820 53618 1876 53630
rect 1820 53566 1822 53618
rect 1874 53566 1876 53618
rect 1820 53172 1876 53566
rect 1820 53078 1876 53116
rect 1820 50484 1876 50494
rect 1820 50034 1876 50428
rect 2044 50372 2100 53788
rect 2156 53506 2212 53518
rect 2156 53454 2158 53506
rect 2210 53454 2212 53506
rect 2156 51492 2212 53454
rect 2268 53060 2324 55020
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 3724 53844 3780 53854
rect 3724 53750 3780 53788
rect 4060 53732 4116 53742
rect 4620 53732 4676 53742
rect 4060 53730 4676 53732
rect 4060 53678 4062 53730
rect 4114 53678 4622 53730
rect 4674 53678 4676 53730
rect 4060 53676 4676 53678
rect 4060 53666 4116 53676
rect 3836 53508 3892 53518
rect 2268 52994 2324 53004
rect 3500 53506 3892 53508
rect 3500 53454 3838 53506
rect 3890 53454 3892 53506
rect 3500 53452 3892 53454
rect 2156 51426 2212 51436
rect 3388 51156 3444 51166
rect 2156 50372 2212 50382
rect 2044 50370 2212 50372
rect 2044 50318 2158 50370
rect 2210 50318 2212 50370
rect 2044 50316 2212 50318
rect 2156 50306 2212 50316
rect 1820 49982 1822 50034
rect 1874 49982 1876 50034
rect 1820 49970 1876 49982
rect 2156 48804 2212 48814
rect 2044 48130 2100 48142
rect 2044 48078 2046 48130
rect 2098 48078 2100 48130
rect 2044 47908 2100 48078
rect 2044 47842 2100 47852
rect 2044 47124 2100 47134
rect 1820 45106 1876 45118
rect 1820 45054 1822 45106
rect 1874 45054 1876 45106
rect 1820 44436 1876 45054
rect 1820 44342 1876 44380
rect 2044 42196 2100 47068
rect 2156 45330 2212 48748
rect 3052 48244 3108 48254
rect 3052 48242 3332 48244
rect 3052 48190 3054 48242
rect 3106 48190 3332 48242
rect 3052 48188 3332 48190
rect 3052 48178 3108 48188
rect 3276 47234 3332 48188
rect 3276 47182 3278 47234
rect 3330 47182 3332 47234
rect 2156 45278 2158 45330
rect 2210 45278 2212 45330
rect 2156 45266 2212 45278
rect 2492 46564 2548 46574
rect 2492 43708 2548 46508
rect 3164 46564 3220 46574
rect 3164 46470 3220 46508
rect 3276 45668 3332 47182
rect 3276 45602 3332 45612
rect 2268 43652 2548 43708
rect 2156 42196 2212 42206
rect 2044 42194 2212 42196
rect 2044 42142 2158 42194
rect 2210 42142 2212 42194
rect 2044 42140 2212 42142
rect 2156 42130 2212 42140
rect 1820 41970 1876 41982
rect 1820 41918 1822 41970
rect 1874 41918 1876 41970
rect 1820 41860 1876 41918
rect 1820 41298 1876 41804
rect 1820 41246 1822 41298
rect 1874 41246 1876 41298
rect 1820 41234 1876 41246
rect 2156 39060 2212 39070
rect 2268 39060 2324 43652
rect 2156 39058 2324 39060
rect 2156 39006 2158 39058
rect 2210 39006 2324 39058
rect 2156 39004 2324 39006
rect 2156 38994 2212 39004
rect 1820 38834 1876 38846
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 38276 1876 38782
rect 1820 38162 1876 38220
rect 1820 38110 1822 38162
rect 1874 38110 1876 38162
rect 1820 38098 1876 38110
rect 1820 36372 1876 36382
rect 1708 36370 1876 36372
rect 1708 36318 1822 36370
rect 1874 36318 1876 36370
rect 1708 36316 1876 36318
rect 1708 35812 1764 36316
rect 1820 36306 1876 36316
rect 1708 35718 1764 35756
rect 2156 36258 2212 36270
rect 2156 36206 2158 36258
rect 2210 36206 2212 36258
rect 2156 34244 2212 36206
rect 3388 35924 3444 51100
rect 3500 36484 3556 53452
rect 3836 53442 3892 53452
rect 3724 53060 3780 53070
rect 3724 52966 3780 53004
rect 3948 53058 4004 53070
rect 3948 53006 3950 53058
rect 4002 53006 4004 53058
rect 3836 52834 3892 52846
rect 3836 52782 3838 52834
rect 3890 52782 3892 52834
rect 3724 51154 3780 51166
rect 3724 51102 3726 51154
rect 3778 51102 3780 51154
rect 3724 48804 3780 51102
rect 3724 48738 3780 48748
rect 3724 48018 3780 48030
rect 3724 47966 3726 48018
rect 3778 47966 3780 48018
rect 3724 47124 3780 47966
rect 3836 47348 3892 52782
rect 3948 52836 4004 53006
rect 3948 51490 4004 52780
rect 3948 51438 3950 51490
rect 4002 51438 4004 51490
rect 3948 50372 4004 51438
rect 3948 50306 4004 50316
rect 4060 51154 4116 51166
rect 4060 51102 4062 51154
rect 4114 51102 4116 51154
rect 4060 49028 4116 51102
rect 4060 48962 4116 48972
rect 4172 48804 4228 53676
rect 4620 53666 4676 53676
rect 6188 53060 6244 53070
rect 6188 52966 6244 53004
rect 4508 52836 4564 52846
rect 4508 52742 4564 52780
rect 5404 52722 5460 52734
rect 5404 52670 5406 52722
rect 5458 52670 5460 52722
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4620 51492 4676 51502
rect 4620 51398 4676 51436
rect 5180 51266 5236 51278
rect 5180 51214 5182 51266
rect 5234 51214 5236 51266
rect 4732 51156 4788 51194
rect 4732 51090 4788 51100
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5180 50372 5236 51214
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4956 49028 5012 49038
rect 4060 48748 4228 48804
rect 4508 48804 4564 48814
rect 3948 48356 4004 48394
rect 3948 48290 4004 48300
rect 3836 47282 3892 47292
rect 3948 48130 4004 48142
rect 3948 48078 3950 48130
rect 4002 48078 4004 48130
rect 3724 47058 3780 47068
rect 3724 46676 3780 46714
rect 3724 46610 3780 46620
rect 3724 46450 3780 46462
rect 3724 46398 3726 46450
rect 3778 46398 3780 46450
rect 3724 43708 3780 46398
rect 3612 43652 3780 43708
rect 3612 36708 3668 43652
rect 3948 39508 4004 48078
rect 4060 46900 4116 48748
rect 4508 48466 4564 48748
rect 4508 48414 4510 48466
rect 4562 48414 4564 48466
rect 4508 48356 4564 48414
rect 4508 48290 4564 48300
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4844 47348 4900 47358
rect 4508 46900 4564 46910
rect 4060 46898 4564 46900
rect 4060 46846 4510 46898
rect 4562 46846 4564 46898
rect 4060 46844 4564 46846
rect 4060 46786 4116 46844
rect 4060 46734 4062 46786
rect 4114 46734 4116 46786
rect 4060 46722 4116 46734
rect 4172 43708 4228 46844
rect 4508 46834 4564 46844
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4172 43652 4340 43708
rect 3948 39442 4004 39452
rect 4172 42644 4228 42654
rect 3836 38724 3892 38734
rect 3612 36642 3668 36652
rect 3724 38668 3836 38724
rect 3500 36418 3556 36428
rect 3388 35858 3444 35868
rect 2156 34178 2212 34188
rect 3500 35476 3556 35486
rect 3500 32788 3556 35420
rect 3052 32786 3556 32788
rect 3052 32734 3502 32786
rect 3554 32734 3556 32786
rect 3052 32732 3556 32734
rect 3052 32562 3108 32732
rect 3500 32722 3556 32732
rect 3052 32510 3054 32562
rect 3106 32510 3108 32562
rect 3052 32498 3108 32510
rect 2044 32452 2100 32462
rect 2044 32358 2100 32396
rect 2268 30884 2324 30894
rect 2156 30324 2212 30334
rect 1820 30098 1876 30110
rect 1820 30046 1822 30098
rect 1874 30046 1876 30098
rect 1820 29652 1876 30046
rect 2156 30098 2212 30268
rect 2156 30046 2158 30098
rect 2210 30046 2212 30098
rect 2156 30034 2212 30046
rect 1820 29558 1876 29596
rect 2156 26962 2212 26974
rect 2156 26910 2158 26962
rect 2210 26910 2212 26962
rect 2156 26404 2212 26910
rect 2156 26338 2212 26348
rect 2156 23826 2212 23838
rect 2156 23774 2158 23826
rect 2210 23774 2212 23826
rect 2156 23716 2212 23774
rect 2156 23650 2212 23660
rect 2044 21474 2100 21486
rect 2044 21422 2046 21474
rect 2098 21422 2100 21474
rect 2044 21028 2100 21422
rect 2044 20962 2100 20972
rect 2156 18676 2212 18686
rect 1820 17556 1876 17566
rect 1820 17106 1876 17500
rect 2156 17554 2212 18620
rect 2156 17502 2158 17554
rect 2210 17502 2212 17554
rect 2156 17490 2212 17502
rect 1820 17054 1822 17106
rect 1874 17054 1876 17106
rect 1820 17042 1876 17054
rect 2156 15540 2212 15550
rect 2268 15540 2324 30828
rect 3500 27188 3556 27198
rect 3724 27188 3780 38668
rect 3836 38592 3892 38668
rect 3948 38612 4004 38622
rect 3948 38518 4004 38556
rect 3836 36708 3892 36718
rect 4172 36708 4228 42588
rect 4284 38164 4340 43652
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4844 39060 4900 47292
rect 4956 39172 5012 48972
rect 5180 48804 5236 50316
rect 5180 48738 5236 48748
rect 5404 47572 5460 52670
rect 7196 52162 7252 56028
rect 7532 56018 7588 56028
rect 12236 56082 12292 56094
rect 12236 56030 12238 56082
rect 12290 56030 12292 56082
rect 7196 52110 7198 52162
rect 7250 52110 7252 52162
rect 6636 48804 6692 48814
rect 6300 48802 6692 48804
rect 6300 48750 6638 48802
rect 6690 48750 6692 48802
rect 6300 48748 6692 48750
rect 5404 47506 5460 47516
rect 5852 47572 5908 47582
rect 5404 44882 5460 44894
rect 5404 44830 5406 44882
rect 5458 44830 5460 44882
rect 5404 43708 5460 44830
rect 5404 43652 5572 43708
rect 5404 43314 5460 43326
rect 5404 43262 5406 43314
rect 5458 43262 5460 43314
rect 4956 39116 5124 39172
rect 4844 38994 4900 39004
rect 4396 38724 4452 38734
rect 4396 38630 4452 38668
rect 5068 38500 5124 39116
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 5068 38434 5124 38444
rect 4476 38378 4740 38388
rect 4284 38108 4900 38164
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4172 36652 4564 36708
rect 3836 36614 3892 36652
rect 4060 36596 4116 36606
rect 4060 36502 4116 36540
rect 4508 36594 4564 36652
rect 4508 36542 4510 36594
rect 4562 36542 4564 36594
rect 4508 36530 4564 36542
rect 4396 36482 4452 36494
rect 4396 36430 4398 36482
rect 4450 36430 4452 36482
rect 4396 36372 4452 36430
rect 4396 36306 4452 36316
rect 4508 36260 4564 36270
rect 4508 36166 4564 36204
rect 4732 36258 4788 36270
rect 4732 36206 4734 36258
rect 4786 36206 4788 36258
rect 4732 36036 4788 36206
rect 4732 35970 4788 35980
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35252 4900 38108
rect 5068 37154 5124 37166
rect 5068 37102 5070 37154
rect 5122 37102 5124 37154
rect 5068 36372 5124 37102
rect 5068 36306 5124 36316
rect 5292 36036 5348 36046
rect 5292 35922 5348 35980
rect 5292 35870 5294 35922
rect 5346 35870 5348 35922
rect 5292 35858 5348 35870
rect 4844 35196 5124 35252
rect 4732 34244 4788 34254
rect 4732 34150 4788 34188
rect 5068 34130 5124 35196
rect 5404 34244 5460 43262
rect 5516 35364 5572 43652
rect 5628 36708 5684 36718
rect 5628 36594 5684 36652
rect 5628 36542 5630 36594
rect 5682 36542 5684 36594
rect 5628 36530 5684 36542
rect 5516 35298 5572 35308
rect 5404 34188 5684 34244
rect 5068 34078 5070 34130
rect 5122 34078 5124 34130
rect 4956 34020 5012 34030
rect 5068 34020 5124 34078
rect 5516 34020 5572 34030
rect 5068 34018 5572 34020
rect 5068 33966 5518 34018
rect 5570 33966 5572 34018
rect 5068 33964 5572 33966
rect 4956 33926 5012 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5516 30996 5572 33964
rect 5628 31892 5684 34188
rect 5628 31826 5684 31836
rect 5516 30930 5572 30940
rect 4732 30884 4788 30894
rect 4732 30790 4788 30828
rect 5180 30884 5236 30894
rect 5180 30790 5236 30828
rect 5516 30770 5572 30782
rect 5516 30718 5518 30770
rect 5570 30718 5572 30770
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5516 30436 5572 30718
rect 5516 30370 5572 30380
rect 5740 30324 5796 30334
rect 5740 30230 5796 30268
rect 5852 30100 5908 47516
rect 6188 45220 6244 45230
rect 6188 45126 6244 45164
rect 6188 43764 6244 43802
rect 6188 43698 6244 43708
rect 6188 40964 6244 40974
rect 5964 30884 6020 30894
rect 5964 30790 6020 30828
rect 5740 30044 5908 30100
rect 5964 30548 6020 30558
rect 5964 30098 6020 30492
rect 6076 30324 6132 30334
rect 6076 30230 6132 30268
rect 5964 30046 5966 30098
rect 6018 30046 6020 30098
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3500 27186 3780 27188
rect 3500 27134 3502 27186
rect 3554 27134 3780 27186
rect 3500 27132 3780 27134
rect 3052 27074 3108 27086
rect 3052 27022 3054 27074
rect 3106 27022 3108 27074
rect 3052 26964 3108 27022
rect 3052 26898 3108 26908
rect 3500 26964 3556 27132
rect 3500 26898 3556 26908
rect 5740 26908 5796 30044
rect 5964 30034 6020 30046
rect 6076 28084 6132 28094
rect 6076 27990 6132 28028
rect 6076 27748 6132 27758
rect 6076 27654 6132 27692
rect 5740 26852 5908 26908
rect 2156 15538 2324 15540
rect 2156 15486 2158 15538
rect 2210 15486 2324 15538
rect 2156 15484 2324 15486
rect 2380 26628 2436 26638
rect 2156 15474 2212 15484
rect 1820 15314 1876 15326
rect 1820 15262 1822 15314
rect 1874 15262 1876 15314
rect 1820 14756 1876 15262
rect 1820 14642 1876 14700
rect 1820 14590 1822 14642
rect 1874 14590 1876 14642
rect 1820 14578 1876 14590
rect 2044 12066 2100 12078
rect 2044 12014 2046 12066
rect 2098 12014 2100 12066
rect 2044 11620 2100 12014
rect 2044 11554 2100 11564
rect 2156 9268 2212 9278
rect 2380 9268 2436 26572
rect 4284 26068 4340 26078
rect 3052 24052 3108 24062
rect 3052 23938 3108 23996
rect 3612 24052 3668 24062
rect 3612 23958 3668 23996
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 3052 23874 3108 23886
rect 3500 23716 3556 23726
rect 3500 21810 3556 23660
rect 3500 21758 3502 21810
rect 3554 21758 3556 21810
rect 3052 21588 3108 21598
rect 3500 21588 3556 21758
rect 3052 21586 3556 21588
rect 3052 21534 3054 21586
rect 3106 21534 3556 21586
rect 3052 21532 3556 21534
rect 3612 22372 3668 22382
rect 3052 21522 3108 21532
rect 3052 12404 3108 12414
rect 3052 12178 3108 12348
rect 3500 12404 3556 12414
rect 3500 12310 3556 12348
rect 3052 12126 3054 12178
rect 3106 12126 3108 12178
rect 3052 12114 3108 12126
rect 2156 9266 2436 9268
rect 2156 9214 2158 9266
rect 2210 9214 2436 9266
rect 2156 9212 2436 9214
rect 2156 9202 2212 9212
rect 1820 9042 1876 9054
rect 1820 8990 1822 9042
rect 1874 8990 1876 9042
rect 1820 8708 1876 8990
rect 1820 8370 1876 8652
rect 3612 8428 3668 22316
rect 3948 21812 4004 21822
rect 3724 20578 3780 20590
rect 3724 20526 3726 20578
rect 3778 20526 3780 20578
rect 3724 18676 3780 20526
rect 3948 20188 4004 21756
rect 4284 20914 4340 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5852 24052 5908 26852
rect 5852 23986 5908 23996
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20862 4286 20914
rect 4338 20862 4340 20914
rect 4284 20850 4340 20862
rect 3948 20132 4340 20188
rect 3724 18610 3780 18620
rect 1820 8318 1822 8370
rect 1874 8318 1876 8370
rect 1820 8306 1876 8318
rect 3388 8372 3668 8428
rect 3052 6132 3108 6142
rect 3052 5906 3108 6076
rect 3052 5854 3054 5906
rect 3106 5854 3108 5906
rect 3052 5842 3108 5854
rect 2044 5794 2100 5806
rect 2044 5742 2046 5794
rect 2098 5742 2100 5794
rect 2044 5572 2100 5742
rect 2044 5506 2100 5516
rect 3052 5236 3108 5246
rect 3052 5122 3108 5180
rect 3052 5070 3054 5122
rect 3106 5070 3108 5122
rect 3052 5058 3108 5070
rect 812 5012 868 5022
rect 140 812 308 868
rect 140 800 196 812
rect -56 728 196 800
rect 252 756 308 812
rect 812 756 868 4956
rect 2156 5012 2212 5022
rect 2156 4918 2212 4956
rect 3388 4564 3444 8372
rect 3500 6132 3556 6142
rect 3500 6038 3556 6076
rect 3612 5236 3668 5246
rect 3612 5142 3668 5180
rect 3500 4564 3556 4574
rect 3388 4562 3556 4564
rect 3388 4510 3502 4562
rect 3554 4510 3556 4562
rect 3388 4508 3556 4510
rect 3052 4340 3108 4350
rect 3388 4340 3444 4508
rect 3500 4498 3556 4508
rect 4284 4564 4340 20132
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 6188 5236 6244 40908
rect 6300 35476 6356 48748
rect 6636 48738 6692 48748
rect 6524 48580 6580 48590
rect 6412 36484 6468 36494
rect 6412 36390 6468 36428
rect 6300 35410 6356 35420
rect 6412 31892 6468 31902
rect 6412 31444 6468 31836
rect 6300 30884 6356 30894
rect 6300 28084 6356 30828
rect 6300 28018 6356 28028
rect 6188 5170 6244 5180
rect 6300 27860 6356 27870
rect 4396 4564 4452 4574
rect 4284 4562 4452 4564
rect 4284 4510 4398 4562
rect 4450 4510 4452 4562
rect 4284 4508 4452 4510
rect 3052 4338 3444 4340
rect 3052 4286 3054 4338
rect 3106 4286 3444 4338
rect 3052 4284 3444 4286
rect 3052 4274 3108 4284
rect 2044 4226 2100 4238
rect 2044 4174 2046 4226
rect 2098 4174 2100 4226
rect 2044 2884 2100 4174
rect 4172 3556 4228 3566
rect 4284 3556 4340 4508
rect 4396 4498 4452 4508
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4172 3554 4340 3556
rect 4172 3502 4174 3554
rect 4226 3502 4340 3554
rect 4172 3500 4340 3502
rect 4172 3490 4228 3500
rect 2044 2818 2100 2828
rect 3276 3442 3332 3454
rect 3276 3390 3278 3442
rect 3330 3390 3332 3442
rect 2828 812 2996 868
rect 2828 800 2884 812
rect -56 200 168 728
rect 252 700 868 756
rect 2632 728 2884 800
rect 2940 756 2996 812
rect 3276 756 3332 3390
rect 5068 3444 5124 3454
rect 5740 3444 5796 3454
rect 5068 3442 5796 3444
rect 5068 3390 5070 3442
rect 5122 3390 5742 3442
rect 5794 3390 5796 3442
rect 5068 3388 5796 3390
rect 5068 3378 5124 3388
rect 2632 200 2856 728
rect 2940 700 3332 756
rect 5292 800 5348 3388
rect 5740 3378 5796 3388
rect 6076 3332 6132 3342
rect 6300 3332 6356 27804
rect 6412 6132 6468 31388
rect 6524 30548 6580 48524
rect 6972 45666 7028 45678
rect 6972 45614 6974 45666
rect 7026 45614 7028 45666
rect 6636 42756 6692 42766
rect 6636 42662 6692 42700
rect 6636 40964 6692 40974
rect 6636 40870 6692 40908
rect 6860 36258 6916 36270
rect 6860 36206 6862 36258
rect 6914 36206 6916 36258
rect 6860 35812 6916 36206
rect 6860 35746 6916 35756
rect 6524 30210 6580 30492
rect 6524 30158 6526 30210
rect 6578 30158 6580 30210
rect 6524 30146 6580 30158
rect 6748 27860 6804 27870
rect 6748 27766 6804 27804
rect 6972 26908 7028 45614
rect 7084 42754 7140 42766
rect 7084 42702 7086 42754
rect 7138 42702 7140 42754
rect 7084 42308 7140 42702
rect 7084 42242 7140 42252
rect 7196 39956 7252 52110
rect 7644 55972 7700 55982
rect 12236 55972 12292 56030
rect 12796 55972 12852 55982
rect 12236 55970 12852 55972
rect 12236 55918 12798 55970
rect 12850 55918 12852 55970
rect 12236 55916 12852 55918
rect 7644 55074 7700 55916
rect 12796 55468 12852 55916
rect 12796 55412 13300 55468
rect 10780 55298 10836 55310
rect 10780 55246 10782 55298
rect 10834 55246 10836 55298
rect 7644 55022 7646 55074
rect 7698 55022 7700 55074
rect 7644 51380 7700 55022
rect 8316 55076 8372 55086
rect 8316 54982 8372 55020
rect 10780 55076 10836 55246
rect 11340 55298 11396 55310
rect 11340 55246 11342 55298
rect 11394 55246 11396 55298
rect 11340 55076 11396 55246
rect 11900 55076 11956 55086
rect 11340 55074 11956 55076
rect 11340 55022 11902 55074
rect 11954 55022 11956 55074
rect 11340 55020 11956 55022
rect 10780 55010 10836 55020
rect 11452 54852 11508 54862
rect 11452 54402 11508 54796
rect 11452 54350 11454 54402
rect 11506 54350 11508 54402
rect 11452 54292 11508 54350
rect 11452 54226 11508 54236
rect 8652 53730 8708 53742
rect 8652 53678 8654 53730
rect 8706 53678 8708 53730
rect 8204 52948 8260 52958
rect 7980 51940 8036 51950
rect 7980 51846 8036 51884
rect 7644 51324 8036 51380
rect 7420 48804 7476 48814
rect 7420 48710 7476 48748
rect 7756 45666 7812 45678
rect 7756 45614 7758 45666
rect 7810 45614 7812 45666
rect 7756 45332 7812 45614
rect 7756 45266 7812 45276
rect 7420 44098 7476 44110
rect 7420 44046 7422 44098
rect 7474 44046 7476 44098
rect 7420 43708 7476 44046
rect 7420 43652 7924 43708
rect 7420 40964 7476 40974
rect 7420 40870 7476 40908
rect 7196 39890 7252 39900
rect 7868 38668 7924 43652
rect 7644 38612 7924 38668
rect 7308 36484 7364 36494
rect 7308 36390 7364 36428
rect 7532 36482 7588 36494
rect 7532 36430 7534 36482
rect 7586 36430 7588 36482
rect 7532 36372 7588 36430
rect 7532 36306 7588 36316
rect 7308 28084 7364 28094
rect 7308 27990 7364 28028
rect 7644 27300 7700 38612
rect 7980 36820 8036 51324
rect 8204 50594 8260 52892
rect 8540 52946 8596 52958
rect 8540 52894 8542 52946
rect 8594 52894 8596 52946
rect 8540 52836 8596 52894
rect 8652 52948 8708 53678
rect 9100 53732 9156 53742
rect 9100 53638 9156 53676
rect 11564 53506 11620 53518
rect 11564 53454 11566 53506
rect 11618 53454 11620 53506
rect 11564 53172 11620 53454
rect 11900 53508 11956 55020
rect 12348 55076 12404 55086
rect 12348 54982 12404 55020
rect 12348 54402 12404 54414
rect 12348 54350 12350 54402
rect 12402 54350 12404 54402
rect 12124 53620 12180 53630
rect 12124 53526 12180 53564
rect 11900 53442 11956 53452
rect 11564 53106 11620 53116
rect 12348 53172 12404 54350
rect 12348 53106 12404 53116
rect 12460 53732 12516 53742
rect 10556 53060 10612 53070
rect 8652 52882 8708 52892
rect 9100 52948 9156 52958
rect 9100 52854 9156 52892
rect 9660 52948 9716 52958
rect 8540 52770 8596 52780
rect 9660 52834 9716 52892
rect 9660 52782 9662 52834
rect 9714 52782 9716 52834
rect 9660 52164 9716 52782
rect 10220 52836 10276 52846
rect 10276 52780 10388 52836
rect 10220 52704 10276 52780
rect 9660 52098 9716 52108
rect 10220 52276 10276 52286
rect 10220 52162 10276 52220
rect 10220 52110 10222 52162
rect 10274 52110 10276 52162
rect 10220 52098 10276 52110
rect 10332 50820 10388 52780
rect 10556 52834 10612 53004
rect 10556 52782 10558 52834
rect 10610 52782 10612 52834
rect 10556 52612 10612 52782
rect 10556 52546 10612 52556
rect 12460 52834 12516 53676
rect 12460 52782 12462 52834
rect 12514 52782 12516 52834
rect 11900 52276 11956 52286
rect 11900 52182 11956 52220
rect 10892 52164 10948 52174
rect 10892 52070 10948 52108
rect 11452 52164 11508 52174
rect 11116 51940 11172 51950
rect 11116 51380 11172 51884
rect 11116 51286 11172 51324
rect 10332 50754 10388 50764
rect 8204 50542 8206 50594
rect 8258 50542 8260 50594
rect 8204 50530 8260 50542
rect 8652 50594 8708 50606
rect 8652 50542 8654 50594
rect 8706 50542 8708 50594
rect 8652 50484 8708 50542
rect 8652 50418 8708 50428
rect 11228 50484 11284 50494
rect 11116 50370 11172 50382
rect 11116 50318 11118 50370
rect 11170 50318 11172 50370
rect 11004 49924 11060 49934
rect 11004 49140 11060 49868
rect 11116 49588 11172 50318
rect 11116 49522 11172 49532
rect 10332 49138 11060 49140
rect 10332 49086 11006 49138
rect 11058 49086 11060 49138
rect 10332 49084 11060 49086
rect 9772 49026 9828 49038
rect 9772 48974 9774 49026
rect 9826 48974 9828 49026
rect 9772 48804 9828 48974
rect 10332 49026 10388 49084
rect 11004 49074 11060 49084
rect 10332 48974 10334 49026
rect 10386 48974 10388 49026
rect 10332 48962 10388 48974
rect 9772 48738 9828 48748
rect 10556 48916 10612 48926
rect 10556 48466 10612 48860
rect 11228 48580 11284 50428
rect 11452 49924 11508 52108
rect 11900 51266 11956 51278
rect 11900 51214 11902 51266
rect 11954 51214 11956 51266
rect 11676 50372 11732 50382
rect 11452 49858 11508 49868
rect 11564 50370 11732 50372
rect 11564 50318 11678 50370
rect 11730 50318 11732 50370
rect 11564 50316 11732 50318
rect 11340 48804 11396 48814
rect 11340 48710 11396 48748
rect 11228 48524 11396 48580
rect 10556 48414 10558 48466
rect 10610 48414 10612 48466
rect 10556 48402 10612 48414
rect 8540 47460 8596 47470
rect 8988 47460 9044 47470
rect 8540 47458 8820 47460
rect 8540 47406 8542 47458
rect 8594 47406 8820 47458
rect 8540 47404 8820 47406
rect 8540 47394 8596 47404
rect 8540 45108 8596 45118
rect 8764 45108 8820 47404
rect 8988 47458 9156 47460
rect 8988 47406 8990 47458
rect 9042 47406 9156 47458
rect 8988 47404 9156 47406
rect 8988 47394 9044 47404
rect 9100 46564 9156 47404
rect 8876 45108 8932 45118
rect 8764 45106 8932 45108
rect 8764 45054 8878 45106
rect 8930 45054 8932 45106
rect 8764 45052 8932 45054
rect 8540 45014 8596 45052
rect 7980 36754 8036 36764
rect 8092 44100 8148 44110
rect 8092 36594 8148 44044
rect 8204 44098 8260 44110
rect 8204 44046 8206 44098
rect 8258 44046 8260 44098
rect 8204 43316 8260 44046
rect 8204 43250 8260 43260
rect 8540 43538 8596 43550
rect 8540 43486 8542 43538
rect 8594 43486 8596 43538
rect 8540 43204 8596 43486
rect 8540 43138 8596 43148
rect 8876 43538 8932 45052
rect 9100 43708 9156 46508
rect 9772 46564 9828 46574
rect 9772 46562 9940 46564
rect 9772 46510 9774 46562
rect 9826 46510 9940 46562
rect 9772 46508 9940 46510
rect 9772 46498 9828 46508
rect 9884 45220 9940 46508
rect 10668 46004 10724 46014
rect 11228 46004 11284 46014
rect 10108 45892 10164 45902
rect 10108 45798 10164 45836
rect 10668 45890 10724 45948
rect 10668 45838 10670 45890
rect 10722 45838 10724 45890
rect 10668 45826 10724 45838
rect 11116 45948 11228 46004
rect 9436 45108 9492 45118
rect 9100 43652 9380 43708
rect 8876 43486 8878 43538
rect 8930 43486 8932 43538
rect 8876 43428 8932 43486
rect 8876 42756 8932 43372
rect 8876 42690 8932 42700
rect 8092 36542 8094 36594
rect 8146 36542 8148 36594
rect 8092 36530 8148 36542
rect 8204 38612 8260 38622
rect 7868 36482 7924 36494
rect 7868 36430 7870 36482
rect 7922 36430 7924 36482
rect 7868 32116 7924 36430
rect 8204 36482 8260 38556
rect 8764 37156 8820 37166
rect 8204 36430 8206 36482
rect 8258 36430 8260 36482
rect 8204 36418 8260 36430
rect 8652 37154 8820 37156
rect 8652 37102 8766 37154
rect 8818 37102 8820 37154
rect 8652 37100 8820 37102
rect 8652 36372 8708 37100
rect 8764 37090 8820 37100
rect 8988 36708 9044 36718
rect 8876 36596 8932 36606
rect 8876 36502 8932 36540
rect 8988 36372 9044 36652
rect 7980 36258 8036 36270
rect 7980 36206 7982 36258
rect 8034 36206 8036 36258
rect 7980 35812 8036 36206
rect 8204 35924 8260 35934
rect 8204 35830 8260 35868
rect 7980 35746 8036 35756
rect 8540 35140 8596 35150
rect 7980 34356 8036 34366
rect 7980 34242 8036 34300
rect 8540 34356 8596 35084
rect 7980 34190 7982 34242
rect 8034 34190 8036 34242
rect 7980 34178 8036 34190
rect 8092 34244 8148 34254
rect 8540 34224 8596 34300
rect 8092 34150 8148 34188
rect 8652 33908 8708 36316
rect 8764 36370 9044 36372
rect 8764 36318 8990 36370
rect 9042 36318 9044 36370
rect 8764 36316 9044 36318
rect 8764 36260 8820 36316
rect 8988 36306 9044 36316
rect 9212 36370 9268 36382
rect 9212 36318 9214 36370
rect 9266 36318 9268 36370
rect 8764 35810 8820 36204
rect 9212 36260 9268 36318
rect 9212 36194 9268 36204
rect 8764 35758 8766 35810
rect 8818 35758 8820 35810
rect 8764 35746 8820 35758
rect 8876 35810 8932 35822
rect 8876 35758 8878 35810
rect 8930 35758 8932 35810
rect 8876 34244 8932 35758
rect 9212 35812 9268 35822
rect 9100 35698 9156 35710
rect 9100 35646 9102 35698
rect 9154 35646 9156 35698
rect 8988 35364 9044 35374
rect 8988 35026 9044 35308
rect 8988 34974 8990 35026
rect 9042 34974 9044 35026
rect 8988 34962 9044 34974
rect 9100 34804 9156 35646
rect 9100 34738 9156 34748
rect 8876 34178 8932 34188
rect 8652 33842 8708 33852
rect 7868 32050 7924 32060
rect 8652 33348 8708 33358
rect 8540 31332 8596 31342
rect 8540 30548 8596 31276
rect 8316 30098 8372 30110
rect 8316 30046 8318 30098
rect 8370 30046 8372 30098
rect 7644 26908 7700 27244
rect 6860 26852 7028 26908
rect 7532 26852 7700 26908
rect 7756 29988 7812 29998
rect 8316 29988 8372 30046
rect 8540 30100 8596 30492
rect 8652 30434 8708 33292
rect 9212 32564 9268 35756
rect 9324 32676 9380 43652
rect 9436 33796 9492 45052
rect 9772 44994 9828 45006
rect 9772 44942 9774 44994
rect 9826 44942 9828 44994
rect 9772 44772 9828 44942
rect 9772 43764 9828 44716
rect 9772 43698 9828 43708
rect 9548 43652 9604 43662
rect 9548 42530 9604 43596
rect 9660 43428 9716 43438
rect 9660 43334 9716 43372
rect 9884 43092 9940 45164
rect 10780 45332 10836 45342
rect 10108 44994 10164 45006
rect 10108 44942 10110 44994
rect 10162 44942 10164 44994
rect 10108 43428 10164 44942
rect 10780 44994 10836 45276
rect 10780 44942 10782 44994
rect 10834 44942 10836 44994
rect 10780 44884 10836 44942
rect 10780 44818 10836 44828
rect 10556 44324 10612 44334
rect 10556 44230 10612 44268
rect 11116 44322 11172 45948
rect 11228 45910 11284 45948
rect 11228 45108 11284 45118
rect 11228 45014 11284 45052
rect 11116 44270 11118 44322
rect 11170 44270 11172 44322
rect 10220 43652 10276 43662
rect 10220 43558 10276 43596
rect 10108 43362 10164 43372
rect 10668 43428 10724 43438
rect 9884 43026 9940 43036
rect 10668 42866 10724 43372
rect 10780 43426 10836 43438
rect 10780 43374 10782 43426
rect 10834 43374 10836 43426
rect 10780 43204 10836 43374
rect 11116 43428 11172 44270
rect 11340 43708 11396 48524
rect 11452 48468 11508 48478
rect 11452 47234 11508 48412
rect 11452 47182 11454 47234
rect 11506 47182 11508 47234
rect 11452 47170 11508 47182
rect 11116 43362 11172 43372
rect 11228 43652 11396 43708
rect 10780 43138 10836 43148
rect 10668 42814 10670 42866
rect 10722 42814 10724 42866
rect 9548 42478 9550 42530
rect 9602 42478 9604 42530
rect 9548 42466 9604 42478
rect 10108 42532 10164 42542
rect 10108 42530 10276 42532
rect 10108 42478 10110 42530
rect 10162 42478 10276 42530
rect 10108 42476 10276 42478
rect 10108 42466 10164 42476
rect 9772 41186 9828 41198
rect 9772 41134 9774 41186
rect 9826 41134 9828 41186
rect 9772 41076 9828 41134
rect 9772 41010 9828 41020
rect 9772 36258 9828 36270
rect 9772 36206 9774 36258
rect 9826 36206 9828 36258
rect 9772 35812 9828 36206
rect 10108 36260 10164 36270
rect 10108 36166 10164 36204
rect 9772 35718 9828 35756
rect 9884 36036 9940 36046
rect 9436 33730 9492 33740
rect 9548 35364 9604 35374
rect 9548 34802 9604 35308
rect 9548 34750 9550 34802
rect 9602 34750 9604 34802
rect 9324 32620 9492 32676
rect 9212 32508 9380 32564
rect 8652 30382 8654 30434
rect 8706 30382 8708 30434
rect 8652 30370 8708 30382
rect 9212 30436 9268 30446
rect 9212 30342 9268 30380
rect 8540 30098 9044 30100
rect 8540 30046 8542 30098
rect 8594 30046 9044 30098
rect 8540 30044 9044 30046
rect 8540 30034 8596 30044
rect 7756 29986 8372 29988
rect 7756 29934 7758 29986
rect 7810 29934 8372 29986
rect 7756 29932 8372 29934
rect 6860 23716 6916 26852
rect 6860 23650 6916 23660
rect 7532 12404 7588 26852
rect 7756 26628 7812 29932
rect 8988 29650 9044 30044
rect 8988 29598 8990 29650
rect 9042 29598 9044 29650
rect 8988 29586 9044 29598
rect 9324 29316 9380 32508
rect 9436 30660 9492 32620
rect 9436 30594 9492 30604
rect 9436 30436 9492 30446
rect 9436 30342 9492 30380
rect 9324 29250 9380 29260
rect 9548 26908 9604 34750
rect 9660 34690 9716 34702
rect 9660 34638 9662 34690
rect 9714 34638 9716 34690
rect 9660 33012 9716 34638
rect 9884 34132 9940 35980
rect 10108 35924 10164 35934
rect 10108 35698 10164 35868
rect 10108 35646 10110 35698
rect 10162 35646 10164 35698
rect 10108 35634 10164 35646
rect 10220 35028 10276 42476
rect 10668 42084 10724 42814
rect 11116 42530 11172 42542
rect 11116 42478 11118 42530
rect 11170 42478 11172 42530
rect 11116 42308 11172 42478
rect 10332 42082 11060 42084
rect 10332 42030 10670 42082
rect 10722 42030 11060 42082
rect 10332 42028 11060 42030
rect 10332 41186 10388 42028
rect 10668 42018 10724 42028
rect 11004 41298 11060 42028
rect 11004 41246 11006 41298
rect 11058 41246 11060 41298
rect 11004 41234 11060 41246
rect 10332 41134 10334 41186
rect 10386 41134 10388 41186
rect 10332 41122 10388 41134
rect 10556 40964 10612 40974
rect 10556 40516 10612 40908
rect 10556 40422 10612 40460
rect 10892 38500 10948 38510
rect 10892 37490 10948 38444
rect 10892 37438 10894 37490
rect 10946 37438 10948 37490
rect 10892 37268 10948 37438
rect 10892 37202 10948 37212
rect 10556 36258 10612 36270
rect 10556 36206 10558 36258
rect 10610 36206 10612 36258
rect 10444 35586 10500 35598
rect 10444 35534 10446 35586
rect 10498 35534 10500 35586
rect 10444 35476 10500 35534
rect 10444 35410 10500 35420
rect 10556 35140 10612 36206
rect 10556 35084 11060 35140
rect 10108 34972 10276 35028
rect 9772 34020 9828 34030
rect 9772 33926 9828 33964
rect 9660 32946 9716 32956
rect 9884 32562 9940 34076
rect 9996 34692 10052 34702
rect 9996 34130 10052 34636
rect 9996 34078 9998 34130
rect 10050 34078 10052 34130
rect 9996 34066 10052 34078
rect 9996 33796 10052 33806
rect 9996 32786 10052 33740
rect 9996 32734 9998 32786
rect 10050 32734 10052 32786
rect 9996 32722 10052 32734
rect 10108 32788 10164 34972
rect 10220 34804 10276 34814
rect 10220 34710 10276 34748
rect 10556 34804 10612 34814
rect 10780 34804 10836 34814
rect 10556 34802 10724 34804
rect 10556 34750 10558 34802
rect 10610 34750 10724 34802
rect 10556 34748 10724 34750
rect 10556 34738 10612 34748
rect 10332 34692 10388 34702
rect 10332 34598 10388 34636
rect 10556 34356 10612 34366
rect 10668 34356 10724 34748
rect 10780 34710 10836 34748
rect 10668 34300 10948 34356
rect 10556 34262 10612 34300
rect 10444 34244 10500 34254
rect 10444 34150 10500 34188
rect 10668 34132 10724 34142
rect 10220 34018 10276 34030
rect 10220 33966 10222 34018
rect 10274 33966 10276 34018
rect 10220 33908 10276 33966
rect 10276 33852 10388 33908
rect 10220 33842 10276 33852
rect 10108 32732 10276 32788
rect 9884 32510 9886 32562
rect 9938 32510 9940 32562
rect 9884 32498 9940 32510
rect 10108 32564 10164 32574
rect 10108 32470 10164 32508
rect 9772 32116 9828 32126
rect 9660 30548 9716 30558
rect 9660 30210 9716 30492
rect 9660 30158 9662 30210
rect 9714 30158 9716 30210
rect 9660 29540 9716 30158
rect 9660 29474 9716 29484
rect 9548 26852 9716 26908
rect 7756 26562 7812 26572
rect 9660 24948 9716 26852
rect 9772 25618 9828 32060
rect 9996 30660 10052 30670
rect 9884 30212 9940 30222
rect 9884 30118 9940 30156
rect 9996 30210 10052 30604
rect 9996 30158 9998 30210
rect 10050 30158 10052 30210
rect 9996 30146 10052 30158
rect 10108 30100 10164 30110
rect 10108 30006 10164 30044
rect 10108 27748 10164 27758
rect 10108 27654 10164 27692
rect 10220 26740 10276 32732
rect 10332 32564 10388 33852
rect 10332 32562 10500 32564
rect 10332 32510 10334 32562
rect 10386 32510 10500 32562
rect 10332 32508 10500 32510
rect 10332 32498 10388 32508
rect 10444 31892 10500 32508
rect 10444 31218 10500 31836
rect 10444 31166 10446 31218
rect 10498 31166 10500 31218
rect 10444 30548 10500 31166
rect 10444 30482 10500 30492
rect 10556 32338 10612 32350
rect 10556 32286 10558 32338
rect 10610 32286 10612 32338
rect 10332 30100 10388 30110
rect 10332 27860 10388 30044
rect 10556 29652 10612 32286
rect 10668 30210 10724 34076
rect 10780 33572 10836 33582
rect 10780 32562 10836 33516
rect 10892 32676 10948 34300
rect 10892 32610 10948 32620
rect 10780 32510 10782 32562
rect 10834 32510 10836 32562
rect 10780 32498 10836 32510
rect 11004 32116 11060 35084
rect 11004 32050 11060 32060
rect 11004 31892 11060 31902
rect 11004 31798 11060 31836
rect 10892 31220 10948 31230
rect 10948 31164 11060 31220
rect 10892 31126 10948 31164
rect 10668 30158 10670 30210
rect 10722 30158 10724 30210
rect 10668 30100 10724 30158
rect 10668 30034 10724 30044
rect 10892 29652 10948 29662
rect 10556 29650 10948 29652
rect 10556 29598 10894 29650
rect 10946 29598 10948 29650
rect 10556 29596 10948 29598
rect 10892 29586 10948 29596
rect 11004 29652 11060 31164
rect 11004 29586 11060 29596
rect 10556 29428 10612 29438
rect 10780 29428 10836 29438
rect 11116 29428 11172 42252
rect 11228 34356 11284 43652
rect 11340 43426 11396 43438
rect 11340 43374 11342 43426
rect 11394 43374 11396 43426
rect 11340 43316 11396 43374
rect 11340 42980 11396 43260
rect 11340 42914 11396 42924
rect 11340 40964 11396 40974
rect 11340 40870 11396 40908
rect 11340 38388 11396 38398
rect 11340 36596 11396 38332
rect 11452 37156 11508 37166
rect 11452 37062 11508 37100
rect 11452 36596 11508 36606
rect 11340 36594 11508 36596
rect 11340 36542 11454 36594
rect 11506 36542 11508 36594
rect 11340 36540 11508 36542
rect 11452 36484 11508 36540
rect 11452 36418 11508 36428
rect 11340 35586 11396 35598
rect 11340 35534 11342 35586
rect 11394 35534 11396 35586
rect 11340 35476 11396 35534
rect 11340 35410 11396 35420
rect 11228 34290 11284 34300
rect 11340 35140 11396 35150
rect 11228 34132 11284 34142
rect 11228 33460 11284 34076
rect 11228 33394 11284 33404
rect 10332 27794 10388 27804
rect 10444 29372 10556 29428
rect 10332 27636 10388 27646
rect 10332 27542 10388 27580
rect 10444 27412 10500 29372
rect 10556 29296 10612 29372
rect 10668 29426 10836 29428
rect 10668 29374 10782 29426
rect 10834 29374 10836 29426
rect 10668 29372 10836 29374
rect 10556 28644 10612 28654
rect 10556 27858 10612 28588
rect 10556 27806 10558 27858
rect 10610 27806 10612 27858
rect 10556 27794 10612 27806
rect 10220 26674 10276 26684
rect 10332 27356 10500 27412
rect 10220 26516 10276 26526
rect 10220 26068 10276 26460
rect 10220 26002 10276 26012
rect 9772 25566 9774 25618
rect 9826 25566 9828 25618
rect 9772 25554 9828 25566
rect 9772 25396 9828 25406
rect 9772 25302 9828 25340
rect 9996 25394 10052 25406
rect 9996 25342 9998 25394
rect 10050 25342 10052 25394
rect 9772 24948 9828 24958
rect 9660 24946 9828 24948
rect 9660 24894 9774 24946
rect 9826 24894 9828 24946
rect 9660 24892 9828 24894
rect 9772 24500 9828 24892
rect 9436 24498 9828 24500
rect 9436 24446 9774 24498
rect 9826 24446 9828 24498
rect 9436 24444 9828 24446
rect 9436 22484 9492 24444
rect 9772 24434 9828 24444
rect 9772 23268 9828 23278
rect 9996 23268 10052 25342
rect 10332 25396 10388 27356
rect 10556 26964 10612 26974
rect 10332 24946 10388 25340
rect 10332 24894 10334 24946
rect 10386 24894 10388 24946
rect 10332 24882 10388 24894
rect 10444 26852 10612 26908
rect 9772 23266 10052 23268
rect 9772 23214 9774 23266
rect 9826 23214 10052 23266
rect 9772 23212 10052 23214
rect 10444 23492 10500 26852
rect 10668 26628 10724 29372
rect 10780 29362 10836 29372
rect 10892 29372 11172 29428
rect 11228 32562 11284 32574
rect 11228 32510 11230 32562
rect 11282 32510 11284 32562
rect 11228 29426 11284 32510
rect 11340 31220 11396 35084
rect 11564 35140 11620 50316
rect 11676 50306 11732 50316
rect 11900 49588 11956 51214
rect 12236 50482 12292 50494
rect 12236 50430 12238 50482
rect 12290 50430 12292 50482
rect 12236 49924 12292 50430
rect 12236 49792 12292 49868
rect 11900 49522 11956 49532
rect 12124 48468 12180 48478
rect 12124 48374 12180 48412
rect 12012 47234 12068 47246
rect 12012 47182 12014 47234
rect 12066 47182 12068 47234
rect 11676 45892 11732 45902
rect 11676 45798 11732 45836
rect 11676 44098 11732 44110
rect 11676 44046 11678 44098
rect 11730 44046 11732 44098
rect 11676 43428 11732 44046
rect 12012 43708 12068 47182
rect 12348 46564 12404 46574
rect 12348 46470 12404 46508
rect 12124 44324 12180 44334
rect 12180 44268 12292 44324
rect 12124 44230 12180 44268
rect 11676 43362 11732 43372
rect 11788 43652 12068 43708
rect 11788 37380 11844 43652
rect 12124 43428 12180 43438
rect 12124 43334 12180 43372
rect 12236 38668 12292 44268
rect 12236 38612 12404 38668
rect 11788 37314 11844 37324
rect 12012 38276 12068 38286
rect 12012 38162 12068 38220
rect 12012 38110 12014 38162
rect 12066 38110 12068 38162
rect 12012 37380 12068 38110
rect 12012 37378 12292 37380
rect 12012 37326 12014 37378
rect 12066 37326 12292 37378
rect 12012 37324 12292 37326
rect 12012 37314 12068 37324
rect 11900 37042 11956 37054
rect 11900 36990 11902 37042
rect 11954 36990 11956 37042
rect 11900 36708 11956 36990
rect 11900 36642 11956 36652
rect 12012 36932 12068 36942
rect 11900 36484 11956 36522
rect 11900 36418 11956 36428
rect 11900 36260 11956 36270
rect 12012 36260 12068 36876
rect 11956 36204 12068 36260
rect 12124 36482 12180 36494
rect 12124 36430 12126 36482
rect 12178 36430 12180 36482
rect 11788 35586 11844 35598
rect 11788 35534 11790 35586
rect 11842 35534 11844 35586
rect 11564 35074 11620 35084
rect 11676 35476 11732 35486
rect 11676 34916 11732 35420
rect 11564 34914 11732 34916
rect 11564 34862 11678 34914
rect 11730 34862 11732 34914
rect 11564 34860 11732 34862
rect 11452 33572 11508 33582
rect 11452 33458 11508 33516
rect 11452 33406 11454 33458
rect 11506 33406 11508 33458
rect 11452 33394 11508 33406
rect 11564 33124 11620 34860
rect 11676 34850 11732 34860
rect 11788 34804 11844 35534
rect 11788 34738 11844 34748
rect 11900 34580 11956 36204
rect 11788 34524 11956 34580
rect 12012 35924 12068 35934
rect 11676 34018 11732 34030
rect 11676 33966 11678 34018
rect 11730 33966 11732 34018
rect 11676 33908 11732 33966
rect 11676 33842 11732 33852
rect 11564 33068 11732 33124
rect 11452 32788 11508 32798
rect 11452 32694 11508 32732
rect 11564 32676 11620 32686
rect 11564 32582 11620 32620
rect 11676 31780 11732 33068
rect 11340 31154 11396 31164
rect 11564 31724 11732 31780
rect 11788 31780 11844 34524
rect 11900 33460 11956 33470
rect 11900 33236 11956 33404
rect 11900 33170 11956 33180
rect 12012 32788 12068 35868
rect 11900 32732 12068 32788
rect 12124 32788 12180 36430
rect 12236 36036 12292 37324
rect 12236 35970 12292 35980
rect 12236 35700 12292 35710
rect 12236 35026 12292 35644
rect 12236 34974 12238 35026
rect 12290 34974 12292 35026
rect 12236 34962 12292 34974
rect 12236 32788 12292 32798
rect 12124 32786 12292 32788
rect 12124 32734 12238 32786
rect 12290 32734 12292 32786
rect 12124 32732 12292 32734
rect 11900 31892 11956 32732
rect 12236 32722 12292 32732
rect 11900 31826 11956 31836
rect 12012 32562 12068 32574
rect 12012 32510 12014 32562
rect 12066 32510 12068 32562
rect 11340 30996 11396 31006
rect 11396 30940 11508 30996
rect 11340 30902 11396 30940
rect 11228 29374 11230 29426
rect 11282 29374 11284 29426
rect 10892 28082 10948 29372
rect 11228 29362 11284 29374
rect 11340 29988 11396 29998
rect 11340 29428 11396 29932
rect 11340 29362 11396 29372
rect 10892 28030 10894 28082
rect 10946 28030 10948 28082
rect 10892 28018 10948 28030
rect 11116 29204 11172 29214
rect 11452 29204 11508 30940
rect 10556 26572 10724 26628
rect 10780 27858 10836 27870
rect 10780 27806 10782 27858
rect 10834 27806 10836 27858
rect 10556 25620 10612 26572
rect 10780 26516 10836 27806
rect 10668 26460 10836 26516
rect 11004 27860 11060 27870
rect 10668 26068 10724 26460
rect 10780 26292 10836 26302
rect 11004 26292 11060 27804
rect 10780 26290 11060 26292
rect 10780 26238 10782 26290
rect 10834 26238 11060 26290
rect 10780 26236 11060 26238
rect 10780 26226 10836 26236
rect 10892 26068 10948 26078
rect 10668 26012 10892 26068
rect 10668 25620 10724 25630
rect 10556 25618 10724 25620
rect 10556 25566 10670 25618
rect 10722 25566 10724 25618
rect 10556 25564 10724 25566
rect 10668 24948 10724 25564
rect 10892 25506 10948 26012
rect 10892 25454 10894 25506
rect 10946 25454 10948 25506
rect 10892 25442 10948 25454
rect 10780 24948 10836 24958
rect 10668 24946 10836 24948
rect 10668 24894 10782 24946
rect 10834 24894 10836 24946
rect 10668 24892 10836 24894
rect 10780 24882 10836 24892
rect 9772 23202 9828 23212
rect 10444 23154 10500 23436
rect 10444 23102 10446 23154
rect 10498 23102 10500 23154
rect 10444 23090 10500 23102
rect 10556 24836 10612 24846
rect 9436 22482 10164 22484
rect 9436 22430 9438 22482
rect 9490 22430 10164 22482
rect 9436 22428 10164 22430
rect 9436 21812 9492 22428
rect 10108 22370 10164 22428
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 22306 10164 22318
rect 10332 22372 10388 22382
rect 10332 22278 10388 22316
rect 10556 22372 10612 24780
rect 10892 24834 10948 24846
rect 10892 24782 10894 24834
rect 10946 24782 10948 24834
rect 10668 24500 10724 24510
rect 10892 24500 10948 24782
rect 11116 24724 11172 29148
rect 11228 29148 11508 29204
rect 11564 29652 11620 31724
rect 11788 31714 11844 31724
rect 11900 31668 11956 31678
rect 11900 31574 11956 31612
rect 11676 31556 11732 31566
rect 11676 30212 11732 31500
rect 11788 31554 11844 31566
rect 11788 31502 11790 31554
rect 11842 31502 11844 31554
rect 11788 30436 11844 31502
rect 12012 31332 12068 32510
rect 12236 32564 12292 32574
rect 11788 30370 11844 30380
rect 11900 31276 12068 31332
rect 12124 31892 12180 31902
rect 11676 30156 11844 30212
rect 11676 29652 11732 29662
rect 11564 29650 11732 29652
rect 11564 29598 11678 29650
rect 11730 29598 11732 29650
rect 11564 29596 11732 29598
rect 11228 24836 11284 29148
rect 11340 28866 11396 28878
rect 11340 28814 11342 28866
rect 11394 28814 11396 28866
rect 11340 28754 11396 28814
rect 11564 28866 11620 29596
rect 11676 29586 11732 29596
rect 11564 28814 11566 28866
rect 11618 28814 11620 28866
rect 11564 28802 11620 28814
rect 11340 28702 11342 28754
rect 11394 28702 11396 28754
rect 11340 28690 11396 28702
rect 11564 27860 11620 27870
rect 11564 27766 11620 27804
rect 11452 27636 11508 27646
rect 11452 27186 11508 27580
rect 11452 27134 11454 27186
rect 11506 27134 11508 27186
rect 11452 27122 11508 27134
rect 11676 27076 11732 27086
rect 11788 27076 11844 30156
rect 11900 28868 11956 31276
rect 12012 31108 12068 31118
rect 12012 31014 12068 31052
rect 12124 31106 12180 31836
rect 12124 31054 12126 31106
rect 12178 31054 12180 31106
rect 12124 30996 12180 31054
rect 12124 30930 12180 30940
rect 12012 30772 12068 30782
rect 12236 30772 12292 32508
rect 12348 32452 12404 38612
rect 12460 36708 12516 52782
rect 12684 53508 12740 53518
rect 12684 52164 12740 53452
rect 12684 52098 12740 52108
rect 13244 52724 13300 55412
rect 13804 53732 13860 53742
rect 13804 53506 13860 53676
rect 13804 53454 13806 53506
rect 13858 53454 13860 53506
rect 13356 52724 13412 52734
rect 13244 52722 13412 52724
rect 13244 52670 13358 52722
rect 13410 52670 13412 52722
rect 13244 52668 13412 52670
rect 12684 50484 12740 50494
rect 12684 50390 12740 50428
rect 12796 48804 12852 48814
rect 12572 47234 12628 47246
rect 12572 47182 12574 47234
rect 12626 47182 12628 47234
rect 12572 46004 12628 47182
rect 12572 45938 12628 45948
rect 12684 43540 12740 43550
rect 12684 43426 12740 43484
rect 12684 43374 12686 43426
rect 12738 43374 12740 43426
rect 12684 42644 12740 43374
rect 12684 42578 12740 42588
rect 12684 38948 12740 38958
rect 12684 37826 12740 38892
rect 12796 38052 12852 48748
rect 13132 48692 13188 48702
rect 13020 43540 13076 43550
rect 12908 43538 13076 43540
rect 12908 43486 13022 43538
rect 13074 43486 13076 43538
rect 12908 43484 13076 43486
rect 12908 43428 12964 43484
rect 13020 43474 13076 43484
rect 12908 42866 12964 43372
rect 12908 42814 12910 42866
rect 12962 42814 12964 42866
rect 12908 42756 12964 42814
rect 12908 42690 12964 42700
rect 13132 38948 13188 48636
rect 13244 40516 13300 52668
rect 13356 52658 13412 52668
rect 13804 48692 13860 53454
rect 13804 48626 13860 48636
rect 14028 47572 14084 59200
rect 16940 59164 17108 59200
rect 17724 55970 17780 59276
rect 19404 59200 19656 59304
rect 22792 59304 23016 59800
rect 22792 59220 23044 59304
rect 23100 59276 23492 59332
rect 23100 59220 23156 59276
rect 22792 59200 23156 59220
rect 19292 56308 19348 56318
rect 19404 56308 19460 59200
rect 22988 59164 23156 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19292 56306 19796 56308
rect 19292 56254 19294 56306
rect 19346 56254 19796 56306
rect 19292 56252 19796 56254
rect 19292 56242 19348 56252
rect 19740 56194 19796 56252
rect 19740 56142 19742 56194
rect 19794 56142 19796 56194
rect 19740 56130 19796 56142
rect 20076 56194 20132 56206
rect 20076 56142 20078 56194
rect 20130 56142 20132 56194
rect 17724 55918 17726 55970
rect 17778 55918 17780 55970
rect 17724 55906 17780 55918
rect 18732 56082 18788 56094
rect 18732 56030 18734 56082
rect 18786 56030 18788 56082
rect 18732 55972 18788 56030
rect 18732 55906 18788 55916
rect 18844 55860 18900 55870
rect 15820 55298 15876 55310
rect 15820 55246 15822 55298
rect 15874 55246 15876 55298
rect 15260 55076 15316 55086
rect 14476 53730 14532 53742
rect 14476 53678 14478 53730
rect 14530 53678 14532 53730
rect 14140 53060 14196 53070
rect 14140 52966 14196 53004
rect 14476 52164 14532 53678
rect 14812 53732 14868 53742
rect 14812 53638 14868 53676
rect 15148 52276 15204 52286
rect 14476 52098 14532 52108
rect 15036 52164 15092 52174
rect 15036 50594 15092 52108
rect 15036 50542 15038 50594
rect 15090 50542 15092 50594
rect 15036 50530 15092 50542
rect 15036 49812 15092 49822
rect 15036 49718 15092 49756
rect 15148 48020 15204 52220
rect 15260 49924 15316 55020
rect 15820 52164 15876 55246
rect 16268 55298 16324 55310
rect 16268 55246 16270 55298
rect 16322 55246 16324 55298
rect 16268 54516 16324 55246
rect 16268 54450 16324 54460
rect 17948 55188 18004 55198
rect 17388 53732 17444 53742
rect 17388 53506 17444 53676
rect 17388 53454 17390 53506
rect 17442 53454 17444 53506
rect 17388 53442 17444 53454
rect 17948 53506 18004 55132
rect 18732 55076 18788 55086
rect 18732 54982 18788 55020
rect 18732 53732 18788 53742
rect 18732 53638 18788 53676
rect 18844 53620 18900 55804
rect 19292 55074 19348 55086
rect 19852 55076 19908 55086
rect 19292 55022 19294 55074
rect 19346 55022 19348 55074
rect 19292 54628 19348 55022
rect 19292 54562 19348 54572
rect 19628 55074 19908 55076
rect 19628 55022 19854 55074
rect 19906 55022 19908 55074
rect 19628 55020 19908 55022
rect 20076 55076 20132 56142
rect 23436 56194 23492 59276
rect 25480 59304 25704 59800
rect 25480 59220 25732 59304
rect 25788 59276 26180 59332
rect 25788 59220 25844 59276
rect 25480 59200 25844 59220
rect 25676 59164 25844 59200
rect 23436 56142 23438 56194
rect 23490 56142 23492 56194
rect 23436 56130 23492 56142
rect 26124 56194 26180 59276
rect 28840 59304 29064 59800
rect 31528 59304 31752 59800
rect 34888 59304 35112 59800
rect 37576 59304 37800 59800
rect 28840 59200 29092 59304
rect 29036 56642 29092 59200
rect 31500 59200 31752 59304
rect 34860 59200 35112 59304
rect 37548 59200 37800 59304
rect 40936 59304 41160 59800
rect 40936 59200 41188 59304
rect 43624 59200 43848 59800
rect 46312 59304 46536 59800
rect 46284 59200 46536 59304
rect 49672 59304 49896 59800
rect 52360 59304 52584 59800
rect 49672 59200 49924 59304
rect 29036 56590 29038 56642
rect 29090 56590 29092 56642
rect 29036 56578 29092 56590
rect 29932 56642 29988 56654
rect 29932 56590 29934 56642
rect 29986 56590 29988 56642
rect 26124 56142 26126 56194
rect 26178 56142 26180 56194
rect 26124 56130 26180 56142
rect 28364 56196 28420 56206
rect 24108 56082 24164 56094
rect 24108 56030 24110 56082
rect 24162 56030 24164 56082
rect 20636 55972 20692 55982
rect 20636 55878 20692 55916
rect 22652 55970 22708 55982
rect 22652 55918 22654 55970
rect 22706 55918 22708 55970
rect 22652 55860 22708 55918
rect 22652 55794 22708 55804
rect 22764 55972 22820 55982
rect 20076 55020 20244 55076
rect 17948 53454 17950 53506
rect 18002 53454 18004 53506
rect 16492 52948 16548 52958
rect 16492 52854 16548 52892
rect 17052 52946 17108 52958
rect 17052 52894 17054 52946
rect 17106 52894 17108 52946
rect 16940 52276 16996 52286
rect 15820 52098 15876 52108
rect 16492 52164 16548 52174
rect 16492 52070 16548 52108
rect 16940 52162 16996 52220
rect 16940 52110 16942 52162
rect 16994 52110 16996 52162
rect 16940 52098 16996 52110
rect 17052 52164 17108 52894
rect 17052 52098 17108 52108
rect 17612 52834 17668 52846
rect 17612 52782 17614 52834
rect 17666 52782 17668 52834
rect 17612 52164 17668 52782
rect 17612 52098 17668 52108
rect 17948 51940 18004 53454
rect 18284 53506 18340 53518
rect 18284 53454 18286 53506
rect 18338 53454 18340 53506
rect 17500 51884 18004 51940
rect 18172 52948 18228 52958
rect 18172 52834 18228 52892
rect 18172 52782 18174 52834
rect 18226 52782 18228 52834
rect 15596 50596 15652 50606
rect 15596 50502 15652 50540
rect 15260 49858 15316 49868
rect 15596 49812 15652 49822
rect 15596 49698 15652 49756
rect 15596 49646 15598 49698
rect 15650 49646 15652 49698
rect 15596 48804 15652 49646
rect 15596 48738 15652 48748
rect 15148 47954 15204 47964
rect 14028 47458 14084 47516
rect 14028 47406 14030 47458
rect 14082 47406 14084 47458
rect 14028 47394 14084 47406
rect 16940 46564 16996 46574
rect 16156 45780 16212 45790
rect 16156 45686 16212 45724
rect 16940 45778 16996 46508
rect 16940 45726 16942 45778
rect 16994 45726 16996 45778
rect 16940 45714 16996 45726
rect 15036 44322 15092 44334
rect 15036 44270 15038 44322
rect 15090 44270 15092 44322
rect 14364 44100 14420 44110
rect 14364 44006 14420 44044
rect 15036 43708 15092 44270
rect 15372 44322 15428 44334
rect 15372 44270 15374 44322
rect 15426 44270 15428 44322
rect 15372 44100 15428 44270
rect 15372 44034 15428 44044
rect 14924 43652 15092 43708
rect 16156 43764 16212 43774
rect 16156 43670 16212 43708
rect 13580 43540 13636 43550
rect 13580 43446 13636 43484
rect 13580 42756 13636 42766
rect 13580 42662 13636 42700
rect 14252 42756 14308 42766
rect 14252 42662 14308 42700
rect 14924 41972 14980 43652
rect 16716 43314 16772 43326
rect 16716 43262 16718 43314
rect 16770 43262 16772 43314
rect 15820 43204 15876 43214
rect 14924 41906 14980 41916
rect 15036 41970 15092 41982
rect 15036 41918 15038 41970
rect 15090 41918 15092 41970
rect 15036 41860 15092 41918
rect 15484 41860 15540 41870
rect 15036 41858 15540 41860
rect 15036 41806 15486 41858
rect 15538 41806 15540 41858
rect 15036 41804 15540 41806
rect 15484 41188 15540 41804
rect 15484 41122 15540 41132
rect 13244 40460 13524 40516
rect 12796 37986 12852 37996
rect 13020 38892 13188 38948
rect 13244 38948 13300 38958
rect 12908 37940 12964 37950
rect 12908 37846 12964 37884
rect 12684 37774 12686 37826
rect 12738 37774 12740 37826
rect 12572 37268 12628 37278
rect 12572 37174 12628 37212
rect 12684 36932 12740 37774
rect 12796 37826 12852 37838
rect 12796 37774 12798 37826
rect 12850 37774 12852 37826
rect 12796 37266 12852 37774
rect 13020 37380 13076 38892
rect 13132 38724 13188 38734
rect 13244 38724 13300 38892
rect 13132 38722 13300 38724
rect 13132 38670 13134 38722
rect 13186 38670 13300 38722
rect 13132 38668 13300 38670
rect 13468 38724 13524 40460
rect 13692 38724 13748 38734
rect 13468 38722 13748 38724
rect 13468 38670 13694 38722
rect 13746 38670 13748 38722
rect 13468 38668 13748 38670
rect 14700 38722 14756 38734
rect 14700 38670 14702 38722
rect 14754 38670 14756 38722
rect 14700 38668 14756 38670
rect 13132 38658 13188 38668
rect 13692 38164 13748 38668
rect 14252 38612 14756 38668
rect 15148 38722 15204 38734
rect 15148 38670 15150 38722
rect 15202 38670 15204 38722
rect 13692 38098 13748 38108
rect 14028 38164 14084 38174
rect 13356 38052 13412 38062
rect 13356 37490 13412 37996
rect 13356 37438 13358 37490
rect 13410 37438 13412 37490
rect 13356 37426 13412 37438
rect 13692 37940 13748 37950
rect 12796 37214 12798 37266
rect 12850 37214 12852 37266
rect 12796 37202 12852 37214
rect 12908 37324 13076 37380
rect 13132 37380 13188 37390
rect 12684 36866 12740 36876
rect 12460 36642 12516 36652
rect 12684 36596 12740 36606
rect 12908 36596 12964 37324
rect 12684 36594 12964 36596
rect 12684 36542 12686 36594
rect 12738 36542 12964 36594
rect 12684 36540 12964 36542
rect 13020 37156 13076 37166
rect 12684 36530 12740 36540
rect 12460 36482 12516 36494
rect 12460 36430 12462 36482
rect 12514 36430 12516 36482
rect 12460 35812 12516 36430
rect 12796 36372 12852 36382
rect 12796 36278 12852 36316
rect 12572 36258 12628 36270
rect 12572 36206 12574 36258
rect 12626 36206 12628 36258
rect 12572 35924 12628 36206
rect 12572 35858 12628 35868
rect 12460 35746 12516 35756
rect 12908 35812 12964 35822
rect 13020 35812 13076 37100
rect 12964 35756 13076 35812
rect 12908 35718 12964 35756
rect 12572 35252 12628 35262
rect 12572 34804 12628 35196
rect 12460 32676 12516 32686
rect 12460 32582 12516 32620
rect 12572 32562 12628 34748
rect 13132 32676 13188 37324
rect 13244 37266 13300 37278
rect 13244 37214 13246 37266
rect 13298 37214 13300 37266
rect 13244 37156 13300 37214
rect 13244 37090 13300 37100
rect 13468 37266 13524 37278
rect 13468 37214 13470 37266
rect 13522 37214 13524 37266
rect 13468 36932 13524 37214
rect 12572 32510 12574 32562
rect 12626 32510 12628 32562
rect 12572 32452 12628 32510
rect 12348 32396 12516 32452
rect 12348 31556 12404 31566
rect 12348 31462 12404 31500
rect 12012 30770 12292 30772
rect 12012 30718 12014 30770
rect 12066 30718 12292 30770
rect 12012 30716 12292 30718
rect 12012 30706 12068 30716
rect 12348 30212 12404 30222
rect 12348 30118 12404 30156
rect 12236 30100 12292 30110
rect 12236 30006 12292 30044
rect 12236 29540 12292 29550
rect 12012 28868 12068 28878
rect 11900 28866 12068 28868
rect 11900 28814 12014 28866
rect 12066 28814 12068 28866
rect 11900 28812 12068 28814
rect 12012 28802 12068 28812
rect 12012 28644 12068 28654
rect 12012 28532 12068 28588
rect 12236 28532 12292 29484
rect 12348 28868 12404 28878
rect 12348 28774 12404 28812
rect 12012 28476 12292 28532
rect 12012 28082 12068 28476
rect 12460 28420 12516 32396
rect 12572 29988 12628 32396
rect 13020 32620 13188 32676
rect 13244 36708 13300 36718
rect 13020 32228 13076 32620
rect 13132 32452 13188 32462
rect 13132 32358 13188 32396
rect 12796 32172 13076 32228
rect 12684 31668 12740 31678
rect 12684 31106 12740 31612
rect 12684 31054 12686 31106
rect 12738 31054 12740 31106
rect 12684 31042 12740 31054
rect 12572 29922 12628 29932
rect 12796 30210 12852 32172
rect 13020 32004 13076 32014
rect 13020 30882 13076 31948
rect 13020 30830 13022 30882
rect 13074 30830 13076 30882
rect 13020 30818 13076 30830
rect 13132 30994 13188 31006
rect 13132 30942 13134 30994
rect 13186 30942 13188 30994
rect 12796 30158 12798 30210
rect 12850 30158 12852 30210
rect 12796 30100 12852 30158
rect 13132 30212 13188 30942
rect 13132 30146 13188 30156
rect 12572 28756 12628 28766
rect 12572 28662 12628 28700
rect 12460 28354 12516 28364
rect 12012 28030 12014 28082
rect 12066 28030 12068 28082
rect 12012 28018 12068 28030
rect 11732 27020 11844 27076
rect 12124 27076 12180 27086
rect 11676 26982 11732 27020
rect 12124 26982 12180 27020
rect 11340 26962 11396 26974
rect 11340 26910 11342 26962
rect 11394 26910 11396 26962
rect 11340 26908 11396 26910
rect 12796 26908 12852 30044
rect 13244 29988 13300 36652
rect 13468 36372 13524 36876
rect 13692 36594 13748 37884
rect 14028 37938 14084 38108
rect 14028 37886 14030 37938
rect 14082 37886 14084 37938
rect 14028 37874 14084 37886
rect 14252 38050 14308 38612
rect 14252 37998 14254 38050
rect 14306 37998 14308 38050
rect 14252 37940 14308 37998
rect 14252 37874 14308 37884
rect 14588 38050 14644 38062
rect 14588 37998 14590 38050
rect 14642 37998 14644 38050
rect 13692 36542 13694 36594
rect 13746 36542 13748 36594
rect 13692 36530 13748 36542
rect 13916 37826 13972 37838
rect 13916 37774 13918 37826
rect 13970 37774 13972 37826
rect 13468 36306 13524 36316
rect 13356 35588 13412 35598
rect 13356 35494 13412 35532
rect 13580 32676 13636 32686
rect 13580 30210 13636 32620
rect 13916 32004 13972 37774
rect 14588 37828 14644 37998
rect 15148 37938 15204 38670
rect 15820 38668 15876 43148
rect 16492 42644 16548 42654
rect 16492 42550 16548 42588
rect 16716 42196 16772 43262
rect 16492 42140 16772 42196
rect 17276 42530 17332 42542
rect 17276 42478 17278 42530
rect 17330 42478 17332 42530
rect 15820 38612 16436 38668
rect 15148 37886 15150 37938
rect 15202 37886 15204 37938
rect 14028 37156 14084 37166
rect 14476 37156 14532 37166
rect 14028 37154 14532 37156
rect 14028 37102 14030 37154
rect 14082 37102 14478 37154
rect 14530 37102 14532 37154
rect 14028 37100 14532 37102
rect 14028 36932 14084 37100
rect 14028 36866 14084 36876
rect 14140 36484 14196 36494
rect 14028 36428 14140 36484
rect 14028 35588 14084 36428
rect 14140 36352 14196 36428
rect 14476 36036 14532 37100
rect 14588 37156 14644 37772
rect 15036 37826 15092 37838
rect 15036 37774 15038 37826
rect 15090 37774 15092 37826
rect 14924 37156 14980 37166
rect 14588 37154 14980 37156
rect 14588 37102 14926 37154
rect 14978 37102 14980 37154
rect 14588 37100 14980 37102
rect 14588 36594 14644 37100
rect 14924 37090 14980 37100
rect 15036 37156 15092 37774
rect 15036 37090 15092 37100
rect 14588 36542 14590 36594
rect 14642 36542 14644 36594
rect 14588 36530 14644 36542
rect 14476 35970 14532 35980
rect 15148 36484 15204 37886
rect 15596 37828 15652 37838
rect 15596 37734 15652 37772
rect 15372 37156 15428 37166
rect 15372 37062 15428 37100
rect 14140 35924 14196 35934
rect 14140 35830 14196 35868
rect 14364 35924 14420 35934
rect 14252 35812 14308 35822
rect 14364 35812 14420 35868
rect 14700 35924 14756 35934
rect 14700 35830 14756 35868
rect 14252 35810 14420 35812
rect 14252 35758 14254 35810
rect 14306 35758 14420 35810
rect 14252 35756 14420 35758
rect 14252 35746 14308 35756
rect 14028 35522 14084 35532
rect 13916 31938 13972 31948
rect 13580 30158 13582 30210
rect 13634 30158 13636 30210
rect 13580 30146 13636 30158
rect 13916 31668 13972 31678
rect 13916 30210 13972 31612
rect 13916 30158 13918 30210
rect 13970 30158 13972 30210
rect 13804 30100 13860 30110
rect 13244 29922 13300 29932
rect 13692 30044 13804 30100
rect 12908 28868 12964 28878
rect 12908 28082 12964 28812
rect 13580 28756 13636 28766
rect 13692 28756 13748 30044
rect 13804 30006 13860 30044
rect 13916 29652 13972 30158
rect 14364 30210 14420 35756
rect 15148 35588 15204 36428
rect 15820 36540 16212 36596
rect 15372 36260 15428 36270
rect 15820 36260 15876 36540
rect 15372 36258 15876 36260
rect 15372 36206 15374 36258
rect 15426 36206 15876 36258
rect 15372 36204 15876 36206
rect 15372 36194 15428 36204
rect 15372 35812 15428 35822
rect 15372 35718 15428 35756
rect 15148 35522 15204 35532
rect 15484 35700 15540 35710
rect 15148 35026 15204 35038
rect 15148 34974 15150 35026
rect 15202 34974 15204 35026
rect 15148 32676 15204 34974
rect 15484 34914 15540 35644
rect 15484 34862 15486 34914
rect 15538 34862 15540 34914
rect 15484 34850 15540 34862
rect 15820 35252 15876 36204
rect 15820 34692 15876 35196
rect 15932 36370 15988 36382
rect 15932 36318 15934 36370
rect 15986 36318 15988 36370
rect 15932 35026 15988 36318
rect 16156 36370 16212 36540
rect 16156 36318 16158 36370
rect 16210 36318 16212 36370
rect 16156 36306 16212 36318
rect 16044 36260 16100 36270
rect 16044 36166 16100 36204
rect 16044 36036 16100 36046
rect 16044 35698 16100 35980
rect 16156 35924 16212 35934
rect 16380 35924 16436 38612
rect 16492 38276 16548 42140
rect 16604 41972 16660 41982
rect 16604 41076 16660 41916
rect 16716 41188 16772 41198
rect 16716 41094 16772 41132
rect 16604 40516 16660 41020
rect 16604 39618 16660 40460
rect 16604 39566 16606 39618
rect 16658 39566 16660 39618
rect 16604 39554 16660 39566
rect 16828 40852 16884 40862
rect 16492 38210 16548 38220
rect 16828 37492 16884 40796
rect 17052 39618 17108 39630
rect 17052 39566 17054 39618
rect 17106 39566 17108 39618
rect 17052 39060 17108 39566
rect 17052 38994 17108 39004
rect 17164 39508 17220 39518
rect 16940 37492 16996 37502
rect 16828 37436 16940 37492
rect 16940 37360 16996 37436
rect 16492 37156 16548 37166
rect 16492 37154 16996 37156
rect 16492 37102 16494 37154
rect 16546 37102 16996 37154
rect 16492 37100 16996 37102
rect 16492 37090 16548 37100
rect 16940 36596 16996 37100
rect 17164 36932 17220 39452
rect 17276 38052 17332 42478
rect 17388 41076 17444 41086
rect 17388 40982 17444 41020
rect 17276 37986 17332 37996
rect 17500 37828 17556 51884
rect 18060 51492 18116 51502
rect 18060 50370 18116 51436
rect 18060 50318 18062 50370
rect 18114 50318 18116 50370
rect 18060 50306 18116 50318
rect 18172 48356 18228 52782
rect 18284 52164 18340 53454
rect 18620 53060 18676 53070
rect 18620 52966 18676 53004
rect 18284 51266 18340 52108
rect 18732 51492 18788 51502
rect 18732 51398 18788 51436
rect 18844 51268 18900 53564
rect 19404 54516 19460 54526
rect 18284 51214 18286 51266
rect 18338 51214 18340 51266
rect 18284 50428 18340 51214
rect 18732 51212 18900 51268
rect 18956 52276 19012 52286
rect 18620 50708 18676 50718
rect 18620 50614 18676 50652
rect 18284 50372 18564 50428
rect 18508 49812 18564 50372
rect 18508 49698 18564 49756
rect 18508 49646 18510 49698
rect 18562 49646 18564 49698
rect 18508 49138 18564 49646
rect 18508 49086 18510 49138
rect 18562 49086 18564 49138
rect 18508 49074 18564 49086
rect 18172 48290 18228 48300
rect 18396 48804 18452 48814
rect 18396 47570 18452 48748
rect 18396 47518 18398 47570
rect 18450 47518 18452 47570
rect 18396 47506 18452 47518
rect 17724 44324 17780 44334
rect 17724 43764 17780 44268
rect 17948 44212 18004 44222
rect 17948 44098 18004 44156
rect 17948 44046 17950 44098
rect 18002 44046 18004 44098
rect 17948 44034 18004 44046
rect 18508 44098 18564 44110
rect 18508 44046 18510 44098
rect 18562 44046 18564 44098
rect 17724 43650 17780 43708
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 17724 43586 17780 43598
rect 17612 42756 17668 42766
rect 17612 38500 17668 42700
rect 18060 42644 18116 42654
rect 18060 42550 18116 42588
rect 18508 38668 18564 44046
rect 18732 43316 18788 51212
rect 18956 51156 19012 52220
rect 19180 51940 19236 51950
rect 18844 51100 19012 51156
rect 19068 51938 19236 51940
rect 19068 51886 19182 51938
rect 19234 51886 19236 51938
rect 19068 51884 19236 51886
rect 18844 50036 18900 51100
rect 19068 50260 19124 51884
rect 19180 51874 19236 51884
rect 19404 50428 19460 54460
rect 19628 54404 19684 55020
rect 19852 55010 19908 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54740 20244 55020
rect 20188 54674 20244 54684
rect 20300 55074 20356 55086
rect 20300 55022 20302 55074
rect 20354 55022 20356 55074
rect 20076 54514 20132 54526
rect 20076 54462 20078 54514
rect 20130 54462 20132 54514
rect 20076 54404 20132 54462
rect 20300 54516 20356 55022
rect 20860 55076 20916 55086
rect 20300 54450 20356 54460
rect 20748 54514 20804 54526
rect 20748 54462 20750 54514
rect 20802 54462 20804 54514
rect 19068 50194 19124 50204
rect 19180 50372 19236 50382
rect 18844 49980 19124 50036
rect 18956 49812 19012 49822
rect 18956 49718 19012 49756
rect 19068 46788 19124 49980
rect 19180 49812 19236 50316
rect 19180 49746 19236 49756
rect 19292 50372 19460 50428
rect 19516 54402 20132 54404
rect 19516 54350 19630 54402
rect 19682 54350 20132 54402
rect 19516 54348 20132 54350
rect 20748 54404 20804 54462
rect 19516 52836 19572 54348
rect 19628 54338 19684 54348
rect 20748 54338 20804 54348
rect 20860 53956 20916 55020
rect 20860 53890 20916 53900
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20524 52946 20580 52958
rect 20524 52894 20526 52946
rect 20578 52894 20580 52946
rect 19516 51378 19572 52780
rect 19964 52836 20020 52846
rect 19964 52742 20020 52780
rect 20524 52836 20580 52894
rect 20524 52274 20580 52780
rect 20524 52222 20526 52274
rect 20578 52222 20580 52274
rect 20524 52210 20580 52222
rect 21084 52946 21140 52958
rect 21084 52894 21086 52946
rect 21138 52894 21140 52946
rect 21084 52052 21140 52894
rect 21532 52276 21588 52286
rect 21532 52182 21588 52220
rect 22092 52164 22148 52174
rect 22652 52164 22708 52174
rect 22092 52162 22260 52164
rect 22092 52110 22094 52162
rect 22146 52110 22260 52162
rect 22092 52108 22260 52110
rect 22092 52098 22148 52108
rect 21084 51986 21140 51996
rect 19964 51940 20020 51950
rect 19516 51326 19518 51378
rect 19570 51326 19572 51378
rect 19516 50372 19572 51326
rect 18956 46732 19124 46788
rect 18844 44100 18900 44110
rect 18844 44006 18900 44044
rect 18732 43260 18900 43316
rect 18732 42532 18788 42542
rect 18620 40516 18676 40526
rect 18620 40422 18676 40460
rect 18508 38612 18676 38668
rect 17612 38444 18004 38500
rect 17500 37772 17668 37828
rect 17612 37604 17668 37772
rect 17164 36866 17220 36876
rect 17500 37548 17668 37604
rect 17388 36596 17444 36606
rect 16940 36594 17220 36596
rect 16940 36542 16942 36594
rect 16994 36542 17220 36594
rect 16940 36540 17220 36542
rect 16940 36530 16996 36540
rect 16156 35922 16436 35924
rect 16156 35870 16158 35922
rect 16210 35870 16436 35922
rect 16156 35868 16436 35870
rect 16492 36372 16548 36382
rect 16156 35858 16212 35868
rect 16492 35812 16548 36316
rect 16044 35646 16046 35698
rect 16098 35646 16100 35698
rect 16044 35364 16100 35646
rect 16268 35700 16324 35710
rect 16268 35606 16324 35644
rect 16492 35698 16548 35756
rect 16492 35646 16494 35698
rect 16546 35646 16548 35698
rect 16492 35634 16548 35646
rect 16716 36260 16772 36270
rect 16716 35698 16772 36204
rect 16716 35646 16718 35698
rect 16770 35646 16772 35698
rect 16716 35634 16772 35646
rect 16828 36258 16884 36270
rect 16828 36206 16830 36258
rect 16882 36206 16884 36258
rect 16828 35700 16884 36206
rect 17164 35922 17220 36540
rect 17164 35870 17166 35922
rect 17218 35870 17220 35922
rect 17164 35858 17220 35870
rect 16828 35634 16884 35644
rect 16940 35700 16996 35710
rect 17388 35700 17444 36540
rect 16940 35698 17444 35700
rect 16940 35646 16942 35698
rect 16994 35646 17444 35698
rect 16940 35644 17444 35646
rect 17500 35924 17556 37548
rect 17724 37492 17780 37502
rect 17724 37380 17780 37436
rect 16940 35634 16996 35644
rect 16044 35298 16100 35308
rect 16716 35476 16772 35486
rect 17164 35476 17220 35486
rect 15932 34974 15934 35026
rect 15986 34974 15988 35026
rect 15932 34962 15988 34974
rect 15820 34626 15876 34636
rect 16156 33348 16212 33358
rect 16716 33348 16772 35420
rect 17052 35474 17220 35476
rect 17052 35422 17166 35474
rect 17218 35422 17220 35474
rect 17052 35420 17220 35422
rect 16940 35364 16996 35374
rect 16940 35026 16996 35308
rect 16940 34974 16942 35026
rect 16994 34974 16996 35026
rect 16940 34962 16996 34974
rect 16156 33346 16772 33348
rect 16156 33294 16158 33346
rect 16210 33294 16718 33346
rect 16770 33294 16772 33346
rect 16156 33292 16772 33294
rect 16156 33282 16212 33292
rect 16716 33282 16772 33292
rect 15148 32610 15204 32620
rect 16044 31892 16100 31902
rect 16044 31444 16100 31836
rect 17052 31892 17108 35420
rect 17164 35410 17220 35420
rect 17276 35252 17332 35262
rect 16604 31668 16660 31678
rect 16604 31574 16660 31612
rect 17052 31666 17108 31836
rect 17164 33460 17220 33470
rect 17164 31890 17220 33404
rect 17276 33458 17332 35196
rect 17276 33406 17278 33458
rect 17330 33406 17332 33458
rect 17276 33394 17332 33406
rect 17164 31838 17166 31890
rect 17218 31838 17220 31890
rect 17164 31826 17220 31838
rect 17500 31890 17556 35868
rect 17612 37378 17780 37380
rect 17612 37326 17726 37378
rect 17778 37326 17780 37378
rect 17612 37324 17780 37326
rect 17612 35140 17668 37324
rect 17724 37314 17780 37324
rect 17836 37042 17892 37054
rect 17836 36990 17838 37042
rect 17890 36990 17892 37042
rect 17724 36932 17780 36942
rect 17724 35924 17780 36876
rect 17836 36484 17892 36990
rect 17948 36708 18004 38444
rect 17948 36642 18004 36652
rect 18172 38052 18228 38062
rect 17892 36428 18004 36484
rect 17836 36418 17892 36428
rect 17836 36260 17892 36270
rect 17836 36166 17892 36204
rect 17836 35924 17892 35934
rect 17724 35922 17892 35924
rect 17724 35870 17838 35922
rect 17890 35870 17892 35922
rect 17724 35868 17892 35870
rect 17836 35700 17892 35868
rect 17836 35634 17892 35644
rect 17836 35364 17892 35374
rect 17612 35084 17780 35140
rect 17612 34914 17668 34926
rect 17612 34862 17614 34914
rect 17666 34862 17668 34914
rect 17612 33460 17668 34862
rect 17612 33394 17668 33404
rect 17724 32676 17780 35084
rect 17500 31838 17502 31890
rect 17554 31838 17556 31890
rect 17052 31614 17054 31666
rect 17106 31614 17108 31666
rect 17052 31602 17108 31614
rect 16828 31554 16884 31566
rect 16828 31502 16830 31554
rect 16882 31502 16884 31554
rect 16044 31378 16100 31388
rect 16380 31444 16436 31454
rect 14364 30158 14366 30210
rect 14418 30158 14420 30210
rect 14364 30100 14420 30158
rect 16044 30212 16100 30222
rect 16044 30118 16100 30156
rect 14364 30034 14420 30044
rect 14924 30100 14980 30110
rect 14924 30006 14980 30044
rect 15484 30100 15540 30110
rect 14140 29652 14196 29662
rect 13916 29650 14196 29652
rect 13916 29598 14142 29650
rect 14194 29598 14196 29650
rect 13916 29596 14196 29598
rect 13916 28868 13972 29596
rect 14140 29586 14196 29596
rect 15484 29316 15540 30044
rect 15484 29250 15540 29260
rect 13916 28802 13972 28812
rect 13636 28700 13748 28756
rect 15820 28756 15876 28766
rect 16380 28756 16436 31388
rect 16828 31444 16884 31502
rect 17500 31444 17556 31838
rect 16828 31388 17556 31444
rect 17612 32620 17780 32676
rect 16828 30212 16884 31388
rect 17500 30548 17556 30558
rect 15820 28754 16436 28756
rect 15820 28702 15822 28754
rect 15874 28702 16382 28754
rect 16434 28702 16436 28754
rect 15820 28700 16436 28702
rect 13580 28624 13636 28700
rect 15820 28690 15876 28700
rect 16380 28690 16436 28700
rect 16604 30156 16884 30212
rect 17052 30324 17108 30334
rect 16604 28866 16660 30156
rect 16828 29986 16884 29998
rect 16828 29934 16830 29986
rect 16882 29934 16884 29986
rect 16828 29876 16884 29934
rect 16828 29810 16884 29820
rect 17052 29650 17108 30268
rect 17164 30212 17220 30222
rect 17164 30118 17220 30156
rect 17052 29598 17054 29650
rect 17106 29598 17108 29650
rect 17052 29586 17108 29598
rect 16604 28814 16606 28866
rect 16658 28814 16660 28866
rect 16604 28644 16660 28814
rect 16940 28756 16996 28766
rect 16940 28662 16996 28700
rect 16604 28578 16660 28588
rect 12908 28030 12910 28082
rect 12962 28030 12964 28082
rect 12908 28018 12964 28030
rect 17500 27188 17556 30492
rect 17612 29650 17668 32620
rect 17724 30324 17780 30334
rect 17724 30230 17780 30268
rect 17836 30212 17892 35308
rect 17948 34914 18004 36428
rect 18060 36260 18116 36270
rect 18060 35364 18116 36204
rect 18060 35298 18116 35308
rect 17948 34862 17950 34914
rect 18002 34862 18004 34914
rect 17948 34850 18004 34862
rect 18172 32228 18228 37996
rect 18508 37826 18564 37838
rect 18508 37774 18510 37826
rect 18562 37774 18564 37826
rect 18508 37380 18564 37774
rect 18396 37324 18564 37380
rect 18284 36372 18340 36382
rect 18396 36372 18452 37324
rect 18340 36316 18452 36372
rect 18508 37154 18564 37166
rect 18508 37102 18510 37154
rect 18562 37102 18564 37154
rect 18508 37044 18564 37102
rect 18284 36278 18340 36316
rect 17948 32172 18228 32228
rect 18284 35812 18340 35822
rect 18284 35364 18340 35756
rect 17948 30548 18004 32172
rect 17948 30482 18004 30492
rect 18060 31668 18116 31678
rect 18060 31554 18116 31612
rect 18060 31502 18062 31554
rect 18114 31502 18116 31554
rect 18060 30436 18116 31502
rect 18060 30370 18116 30380
rect 17836 30146 17892 30156
rect 17948 30210 18004 30222
rect 17948 30158 17950 30210
rect 18002 30158 18004 30210
rect 17612 29598 17614 29650
rect 17666 29598 17668 29650
rect 17612 28756 17668 29598
rect 17948 28868 18004 30158
rect 18284 30210 18340 35308
rect 18508 35252 18564 36988
rect 18620 35364 18676 38612
rect 18732 37044 18788 42476
rect 18844 37268 18900 43260
rect 18956 43204 19012 46732
rect 19292 46564 19348 50372
rect 19516 50306 19572 50316
rect 19628 51938 20020 51940
rect 19628 51886 19966 51938
rect 20018 51886 20020 51938
rect 19628 51884 20020 51886
rect 19628 50036 19684 51884
rect 19964 51874 20020 51884
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19740 51604 19796 51614
rect 19740 50596 19796 51548
rect 19740 50502 19796 50540
rect 20188 51378 20244 51390
rect 20188 51326 20190 51378
rect 20242 51326 20244 51378
rect 20188 50372 20244 51326
rect 20188 50306 20244 50316
rect 22092 50932 22148 50942
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19628 49980 19796 50036
rect 19628 49810 19684 49822
rect 19628 49758 19630 49810
rect 19682 49758 19684 49810
rect 19628 49700 19684 49758
rect 19628 49634 19684 49644
rect 19740 48804 19796 49980
rect 22092 50034 22148 50876
rect 22092 49982 22094 50034
rect 22146 49982 22148 50034
rect 22092 49970 22148 49982
rect 22204 50036 22260 52108
rect 22652 51602 22708 52108
rect 22652 51550 22654 51602
rect 22706 51550 22708 51602
rect 22652 51538 22708 51550
rect 22764 50428 22820 55916
rect 24108 55860 24164 56030
rect 24108 55794 24164 55804
rect 25340 56084 25396 56094
rect 23212 54738 23268 54750
rect 23212 54686 23214 54738
rect 23266 54686 23268 54738
rect 23212 53620 23268 54686
rect 24220 54404 24276 54414
rect 24220 54310 24276 54348
rect 23772 54292 23828 54302
rect 23772 54290 24052 54292
rect 23772 54238 23774 54290
rect 23826 54238 24052 54290
rect 23772 54236 24052 54238
rect 23772 54226 23828 54236
rect 23212 53554 23268 53564
rect 23436 53172 23492 53182
rect 23436 53078 23492 53116
rect 23660 51266 23716 51278
rect 23660 51214 23662 51266
rect 23714 51214 23716 51266
rect 19628 48748 19796 48804
rect 20524 49026 20580 49038
rect 20524 48974 20526 49026
rect 20578 48974 20580 49026
rect 20524 48804 20580 48974
rect 19404 47572 19460 47582
rect 19404 47478 19460 47516
rect 19628 46900 19684 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 46844 19796 46900
rect 19292 46508 19572 46564
rect 19180 45892 19236 45902
rect 19180 45798 19236 45836
rect 19404 45668 19460 45678
rect 19292 44212 19348 44222
rect 19292 44118 19348 44156
rect 18956 43148 19236 43204
rect 18956 40964 19012 40974
rect 18956 37492 19012 40908
rect 19068 40516 19124 40526
rect 19068 40402 19124 40460
rect 19068 40350 19070 40402
rect 19122 40350 19124 40402
rect 19068 40338 19124 40350
rect 18956 37426 19012 37436
rect 19068 37826 19124 37838
rect 19068 37774 19070 37826
rect 19122 37774 19124 37826
rect 18844 37202 18900 37212
rect 19068 37044 19124 37774
rect 18732 36978 18788 36988
rect 18844 37042 19124 37044
rect 18844 36990 19070 37042
rect 19122 36990 19124 37042
rect 18844 36988 19124 36990
rect 18732 36260 18788 36270
rect 18732 35922 18788 36204
rect 18732 35870 18734 35922
rect 18786 35870 18788 35922
rect 18732 35858 18788 35870
rect 18620 35308 18788 35364
rect 18508 35196 18676 35252
rect 18508 34804 18564 34814
rect 18508 34710 18564 34748
rect 18620 33236 18676 35196
rect 18620 33170 18676 33180
rect 18284 30158 18286 30210
rect 18338 30158 18340 30210
rect 18284 29876 18340 30158
rect 18620 30212 18676 30222
rect 18620 30118 18676 30156
rect 18284 29810 18340 29820
rect 18396 29986 18452 29998
rect 18396 29934 18398 29986
rect 18450 29934 18452 29986
rect 18396 29652 18452 29934
rect 18508 29988 18564 29998
rect 18508 29894 18564 29932
rect 18732 29764 18788 35308
rect 18844 33348 18900 36988
rect 19068 36978 19124 36988
rect 19180 36708 19236 43148
rect 19292 37492 19348 37502
rect 19292 37266 19348 37436
rect 19404 37380 19460 45612
rect 19516 40292 19572 46508
rect 19628 46562 19684 46574
rect 19628 46510 19630 46562
rect 19682 46510 19684 46562
rect 19628 45890 19684 46510
rect 19628 45838 19630 45890
rect 19682 45838 19684 45890
rect 19628 44996 19684 45838
rect 19740 45668 19796 46844
rect 20412 46674 20468 46686
rect 20412 46622 20414 46674
rect 20466 46622 20468 46674
rect 20076 46564 20132 46574
rect 20076 46470 20132 46508
rect 19740 45602 19796 45612
rect 20412 45666 20468 46622
rect 20412 45614 20414 45666
rect 20466 45614 20468 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45108 20244 45118
rect 20412 45108 20468 45614
rect 20188 45106 20468 45108
rect 20188 45054 20190 45106
rect 20242 45054 20468 45106
rect 20188 45052 20468 45054
rect 19740 44996 19796 45006
rect 20188 44996 20244 45052
rect 19628 44994 20244 44996
rect 19628 44942 19742 44994
rect 19794 44942 20244 44994
rect 19628 44940 20244 44942
rect 19628 44100 19684 44940
rect 19740 44930 19796 44940
rect 19628 43428 19684 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20300 43538 20356 43550
rect 20300 43486 20302 43538
rect 20354 43486 20356 43538
rect 19852 43428 19908 43438
rect 20300 43428 20356 43486
rect 19628 43426 20356 43428
rect 19628 43374 19854 43426
rect 19906 43374 20356 43426
rect 19628 43372 20356 43374
rect 19628 41860 19684 43372
rect 19852 43362 19908 43372
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20076 41970 20132 41982
rect 20076 41918 20078 41970
rect 20130 41918 20132 41970
rect 20076 41860 20132 41918
rect 19628 41858 20132 41860
rect 19628 41806 19630 41858
rect 19682 41806 20132 41858
rect 19628 41804 20132 41806
rect 19628 40516 19684 41804
rect 20524 41188 20580 48748
rect 21532 48804 21588 48814
rect 21532 48710 21588 48748
rect 22204 48804 22260 49980
rect 22204 48738 22260 48748
rect 22652 50372 22820 50428
rect 23212 51154 23268 51166
rect 23212 51102 23214 51154
rect 23266 51102 23268 51154
rect 22652 49586 22708 50372
rect 23100 49700 23156 49710
rect 23100 49606 23156 49644
rect 22652 49534 22654 49586
rect 22706 49534 22708 49586
rect 21084 46674 21140 46686
rect 21084 46622 21086 46674
rect 21138 46622 21140 46674
rect 21084 46452 21140 46622
rect 21084 46386 21140 46396
rect 21868 46004 21924 46014
rect 20860 45892 20916 45902
rect 20860 45666 20916 45836
rect 20860 45614 20862 45666
rect 20914 45614 20916 45666
rect 20748 45108 20804 45118
rect 20748 45014 20804 45052
rect 20524 41122 20580 41132
rect 20748 41970 20804 41982
rect 20748 41918 20750 41970
rect 20802 41918 20804 41970
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40450 19684 40460
rect 20636 40516 20692 40526
rect 19740 40402 19796 40414
rect 19740 40350 19742 40402
rect 19794 40350 19796 40402
rect 19740 40292 19796 40350
rect 19516 40236 19684 40292
rect 19516 39620 19572 39630
rect 19516 39394 19572 39564
rect 19516 39342 19518 39394
rect 19570 39342 19572 39394
rect 19516 39330 19572 39342
rect 19628 37492 19684 40236
rect 19740 40226 19796 40236
rect 20076 39844 20132 39854
rect 20076 39750 20132 39788
rect 20636 39730 20692 40460
rect 20748 40180 20804 41918
rect 20748 40114 20804 40124
rect 20636 39678 20638 39730
rect 20690 39678 20692 39730
rect 20636 39666 20692 39678
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20412 39060 20468 39070
rect 20412 38966 20468 39004
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19852 37492 19908 37502
rect 19628 37490 19908 37492
rect 19628 37438 19854 37490
rect 19906 37438 19908 37490
rect 19628 37436 19908 37438
rect 19852 37426 19908 37436
rect 20524 37492 20580 37502
rect 20524 37398 20580 37436
rect 19404 37324 19684 37380
rect 19292 37214 19294 37266
rect 19346 37214 19348 37266
rect 19292 37202 19348 37214
rect 19516 37156 19572 37166
rect 19404 37154 19572 37156
rect 19404 37102 19518 37154
rect 19570 37102 19572 37154
rect 19404 37100 19572 37102
rect 19180 36652 19348 36708
rect 19068 36596 19124 36606
rect 19068 36502 19124 36540
rect 19180 36484 19236 36494
rect 19180 36390 19236 36428
rect 18956 36260 19012 36270
rect 18956 36166 19012 36204
rect 19180 36148 19236 36158
rect 19068 34804 19124 34814
rect 19068 34710 19124 34748
rect 19180 33348 19236 36092
rect 19292 35924 19348 36652
rect 19404 36484 19460 37100
rect 19516 37090 19572 37100
rect 19628 36932 19684 37324
rect 19740 37268 19796 37278
rect 19740 37174 19796 37212
rect 19964 37266 20020 37278
rect 19964 37214 19966 37266
rect 20018 37214 20020 37266
rect 19964 37044 20020 37214
rect 19964 36978 20020 36988
rect 19404 36390 19460 36428
rect 19516 36876 19684 36932
rect 19516 36260 19572 36876
rect 19852 36596 19908 36606
rect 19852 36502 19908 36540
rect 20412 36596 20468 36606
rect 20412 36502 20468 36540
rect 19292 35858 19348 35868
rect 19404 36204 19572 36260
rect 19628 36482 19684 36494
rect 19628 36430 19630 36482
rect 19682 36430 19684 36482
rect 19292 35700 19348 35710
rect 19292 35606 19348 35644
rect 19404 35364 19460 36204
rect 19292 35308 19460 35364
rect 19516 35474 19572 35486
rect 19516 35422 19518 35474
rect 19570 35422 19572 35474
rect 19516 35364 19572 35422
rect 19292 34916 19348 35308
rect 19516 35298 19572 35308
rect 19404 35140 19460 35150
rect 19628 35140 19684 36430
rect 20188 36260 20244 36270
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20076 35924 20132 35934
rect 20076 35830 20132 35868
rect 19852 35812 19908 35822
rect 19852 35698 19908 35756
rect 19852 35646 19854 35698
rect 19906 35646 19908 35698
rect 19852 35634 19908 35646
rect 19964 35698 20020 35710
rect 19964 35646 19966 35698
rect 20018 35646 20020 35698
rect 19404 35138 19684 35140
rect 19404 35086 19406 35138
rect 19458 35086 19684 35138
rect 19404 35084 19684 35086
rect 19964 35140 20020 35646
rect 20188 35698 20244 36204
rect 20188 35646 20190 35698
rect 20242 35646 20244 35698
rect 20188 35252 20244 35646
rect 20860 35252 20916 45614
rect 20972 43652 21028 43662
rect 20972 43538 21028 43596
rect 20972 43486 20974 43538
rect 21026 43486 21028 43538
rect 20972 43474 21028 43486
rect 21532 41188 21588 41198
rect 21532 41094 21588 41132
rect 21532 39620 21588 39630
rect 21532 39526 21588 39564
rect 21756 39060 21812 39070
rect 20972 37268 21028 37278
rect 20972 37174 21028 37212
rect 21756 35924 21812 39004
rect 21756 35858 21812 35868
rect 20188 35196 20580 35252
rect 20860 35196 21028 35252
rect 19964 35084 20244 35140
rect 19404 35074 19460 35084
rect 19292 34860 19460 34916
rect 19292 34692 19348 34702
rect 19292 34598 19348 34636
rect 19404 34020 19460 34860
rect 19852 34692 19908 34730
rect 19852 34626 19908 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19404 33954 19460 33964
rect 19852 34020 19908 34030
rect 19852 33926 19908 33964
rect 19964 33908 20020 33918
rect 19964 33814 20020 33852
rect 20188 33908 20244 35084
rect 20412 34916 20468 34926
rect 20412 34692 20468 34860
rect 20188 33842 20244 33852
rect 20300 34690 20468 34692
rect 20300 34638 20414 34690
rect 20466 34638 20468 34690
rect 20300 34636 20468 34638
rect 20300 33684 20356 34636
rect 20412 34626 20468 34636
rect 20524 34244 20580 35196
rect 20860 34692 20916 34702
rect 20860 34598 20916 34636
rect 20524 34178 20580 34188
rect 20412 34020 20468 34030
rect 20468 33964 20580 34020
rect 20412 33888 20468 33964
rect 20300 33618 20356 33628
rect 19180 33292 19460 33348
rect 18844 33282 18900 33292
rect 19292 33124 19348 33134
rect 19068 30882 19124 30894
rect 19068 30830 19070 30882
rect 19122 30830 19124 30882
rect 18396 29586 18452 29596
rect 18620 29708 18788 29764
rect 18956 30100 19012 30110
rect 18284 29540 18340 29550
rect 18172 29316 18228 29326
rect 17948 28802 18004 28812
rect 18060 29314 18228 29316
rect 18060 29262 18174 29314
rect 18226 29262 18228 29314
rect 18060 29260 18228 29262
rect 18060 28868 18116 29260
rect 18172 29250 18228 29260
rect 18284 28980 18340 29484
rect 18508 29426 18564 29438
rect 18508 29374 18510 29426
rect 18562 29374 18564 29426
rect 18284 28924 18452 28980
rect 18060 28812 18340 28868
rect 17724 28756 17780 28766
rect 17612 28754 17892 28756
rect 17612 28702 17726 28754
rect 17778 28702 17892 28754
rect 17612 28700 17892 28702
rect 17724 28690 17780 28700
rect 17836 28644 17892 28700
rect 18060 28644 18116 28812
rect 17836 28588 18116 28644
rect 18172 28644 18228 28654
rect 18172 28550 18228 28588
rect 18284 28642 18340 28812
rect 18284 28590 18286 28642
rect 18338 28590 18340 28642
rect 18284 28578 18340 28590
rect 17724 28532 17780 28542
rect 18396 28532 18452 28924
rect 18508 28756 18564 29374
rect 18508 28690 18564 28700
rect 18508 28532 18564 28542
rect 18396 28530 18564 28532
rect 18396 28478 18510 28530
rect 18562 28478 18564 28530
rect 18396 28476 18564 28478
rect 17724 28082 17780 28476
rect 18508 28466 18564 28476
rect 17724 28030 17726 28082
rect 17778 28030 17780 28082
rect 17724 28018 17780 28030
rect 17836 27188 17892 27198
rect 17500 27186 17892 27188
rect 17500 27134 17838 27186
rect 17890 27134 17892 27186
rect 17500 27132 17892 27134
rect 17388 27076 17444 27086
rect 17388 26982 17444 27020
rect 11340 26852 11508 26908
rect 11340 26628 11396 26638
rect 11340 26514 11396 26572
rect 11340 26462 11342 26514
rect 11394 26462 11396 26514
rect 11340 26450 11396 26462
rect 11452 25620 11508 26852
rect 12348 26852 12852 26908
rect 17836 26964 17892 27132
rect 18284 27188 18340 27198
rect 18284 27094 18340 27132
rect 17836 26898 17892 26908
rect 12012 26740 12068 26750
rect 12012 26402 12068 26684
rect 12012 26350 12014 26402
rect 12066 26350 12068 26402
rect 11900 26068 11956 26078
rect 11900 25974 11956 26012
rect 11564 25620 11620 25630
rect 11452 25618 11620 25620
rect 11452 25566 11566 25618
rect 11618 25566 11620 25618
rect 11452 25564 11620 25566
rect 11564 25554 11620 25564
rect 11340 24836 11396 24846
rect 11228 24780 11340 24836
rect 11340 24704 11396 24780
rect 11788 24724 11844 24734
rect 11116 24630 11172 24668
rect 10668 24498 10948 24500
rect 10668 24446 10670 24498
rect 10722 24446 10948 24498
rect 10668 24444 10948 24446
rect 11788 24610 11844 24668
rect 11788 24558 11790 24610
rect 11842 24558 11844 24610
rect 10668 24434 10724 24444
rect 11340 23492 11396 23502
rect 11340 23378 11396 23436
rect 11340 23326 11342 23378
rect 11394 23326 11396 23378
rect 11340 23314 11396 23326
rect 10668 23044 10724 23054
rect 10668 22950 10724 22988
rect 11004 23044 11060 23054
rect 11004 22594 11060 22988
rect 11676 23044 11732 23054
rect 11676 22950 11732 22988
rect 11788 22820 11844 24558
rect 11004 22542 11006 22594
rect 11058 22542 11060 22594
rect 11004 22530 11060 22542
rect 11676 22764 11844 22820
rect 11676 22372 11732 22764
rect 12012 22596 12068 26350
rect 12236 24836 12292 24846
rect 12236 24742 12292 24780
rect 10556 22370 11396 22372
rect 10556 22318 10558 22370
rect 10610 22318 11396 22370
rect 10556 22316 11396 22318
rect 10556 22306 10612 22316
rect 9996 22260 10052 22270
rect 9996 22166 10052 22204
rect 9436 21746 9492 21756
rect 11340 21810 11396 22316
rect 11676 22306 11732 22316
rect 11788 22540 12068 22596
rect 11788 22482 11844 22540
rect 11788 22430 11790 22482
rect 11842 22430 11844 22482
rect 11340 21758 11342 21810
rect 11394 21758 11396 21810
rect 7532 12338 7588 12348
rect 6412 6066 6468 6076
rect 11340 5348 11396 21758
rect 11340 5282 11396 5292
rect 11788 22260 11844 22430
rect 12236 22372 12292 22382
rect 12236 22278 12292 22316
rect 11116 4564 11172 4574
rect 10892 3556 10948 3566
rect 11116 3556 11172 4508
rect 11788 3668 11844 22204
rect 12348 4564 12404 26852
rect 12460 26740 12516 26750
rect 12460 26514 12516 26684
rect 12460 26462 12462 26514
rect 12514 26462 12516 26514
rect 12460 26450 12516 26462
rect 18172 24836 18228 24846
rect 18060 24612 18116 24622
rect 17164 23938 17220 23950
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 17164 23492 17220 23886
rect 17164 23426 17220 23436
rect 17388 23938 17444 23950
rect 17388 23886 17390 23938
rect 17442 23886 17444 23938
rect 17388 23380 17444 23886
rect 17724 23828 17780 23838
rect 17724 23734 17780 23772
rect 17948 23492 18004 23502
rect 17388 23314 17444 23324
rect 17836 23380 17892 23390
rect 17836 23154 17892 23324
rect 17948 23266 18004 23436
rect 18060 23378 18116 24556
rect 18060 23326 18062 23378
rect 18114 23326 18116 23378
rect 18060 23314 18116 23326
rect 18172 24050 18228 24780
rect 18172 23998 18174 24050
rect 18226 23998 18228 24050
rect 18172 23380 18228 23998
rect 18620 24050 18676 29708
rect 18956 29426 19012 30044
rect 19068 29652 19124 30830
rect 19180 30436 19236 30446
rect 19180 30342 19236 30380
rect 19068 29586 19124 29596
rect 19180 29652 19236 29662
rect 19292 29652 19348 33068
rect 19180 29650 19348 29652
rect 19180 29598 19182 29650
rect 19234 29598 19348 29650
rect 19180 29596 19348 29598
rect 19180 29586 19236 29596
rect 19404 29428 19460 33292
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19852 30268 20132 30324
rect 19628 30212 19684 30222
rect 19628 30118 19684 30156
rect 19852 30210 19908 30268
rect 19852 30158 19854 30210
rect 19906 30158 19908 30210
rect 19852 30146 19908 30158
rect 19964 30100 20020 30110
rect 19964 30006 20020 30044
rect 20076 29988 20132 30268
rect 20188 30212 20244 30222
rect 20188 30210 20468 30212
rect 20188 30158 20190 30210
rect 20242 30158 20468 30210
rect 20188 30156 20468 30158
rect 20188 30146 20244 30156
rect 20412 30100 20468 30156
rect 20412 30034 20468 30044
rect 20076 29932 20356 29988
rect 20300 29876 20356 29932
rect 20412 29876 20468 29886
rect 19836 29820 20100 29830
rect 20300 29820 20412 29876
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20412 29650 20468 29820
rect 20412 29598 20414 29650
rect 20466 29598 20468 29650
rect 20412 29586 20468 29598
rect 18956 29374 18958 29426
rect 19010 29374 19012 29426
rect 18732 28756 18788 28766
rect 18732 28642 18788 28700
rect 18956 28644 19012 29374
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 18732 28578 18788 28590
rect 18844 28642 19012 28644
rect 18844 28590 18958 28642
rect 19010 28590 19012 28642
rect 18844 28588 19012 28590
rect 18732 27300 18788 27310
rect 18844 27300 18900 28588
rect 18956 28578 19012 28588
rect 19180 29372 19460 29428
rect 19516 29540 19572 29550
rect 18732 27298 18900 27300
rect 18732 27246 18734 27298
rect 18786 27246 18900 27298
rect 18732 27244 18900 27246
rect 18732 27234 18788 27244
rect 19180 27188 19236 29372
rect 19404 28756 19460 28766
rect 19516 28756 19572 29484
rect 19404 28754 19572 28756
rect 19404 28702 19406 28754
rect 19458 28702 19572 28754
rect 19404 28700 19572 28702
rect 19404 28690 19460 28700
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27860 19572 27870
rect 19180 27074 19236 27132
rect 19180 27022 19182 27074
rect 19234 27022 19236 27074
rect 19180 27010 19236 27022
rect 19404 27188 19460 27198
rect 19404 27074 19460 27132
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 27010 19460 27022
rect 19516 26964 19572 27804
rect 20188 27748 20244 27758
rect 20188 27188 20244 27692
rect 20524 27748 20580 33964
rect 20972 31780 21028 35196
rect 21868 35026 21924 45948
rect 22204 40628 22260 40638
rect 22204 40534 22260 40572
rect 22652 38668 22708 49534
rect 23212 48132 23268 51102
rect 23660 50372 23716 51214
rect 23660 49812 23716 50316
rect 23660 49746 23716 49756
rect 23212 48066 23268 48076
rect 23436 47236 23492 47246
rect 23324 47124 23380 47134
rect 23324 45330 23380 47068
rect 23436 46898 23492 47180
rect 23436 46846 23438 46898
rect 23490 46846 23492 46898
rect 23436 46834 23492 46846
rect 23324 45278 23326 45330
rect 23378 45278 23380 45330
rect 23324 45266 23380 45278
rect 23548 46452 23604 46462
rect 23436 43764 23492 43774
rect 23436 43670 23492 43708
rect 23212 42196 23268 42206
rect 23212 42102 23268 42140
rect 22764 41188 22820 41198
rect 22764 40626 22820 41132
rect 22764 40574 22766 40626
rect 22818 40574 22820 40626
rect 22764 40562 22820 40574
rect 23212 40402 23268 40414
rect 23212 40350 23214 40402
rect 23266 40350 23268 40402
rect 23212 40292 23268 40350
rect 23212 38836 23268 40236
rect 23212 38770 23268 38780
rect 22652 38612 22820 38668
rect 22540 35252 22596 35262
rect 21868 34974 21870 35026
rect 21922 34974 21924 35026
rect 21868 34962 21924 34974
rect 22428 35028 22484 35038
rect 22428 34934 22484 34972
rect 22092 34916 22148 34926
rect 22092 34822 22148 34860
rect 21756 34690 21812 34702
rect 21756 34638 21758 34690
rect 21810 34638 21812 34690
rect 21756 34580 21812 34638
rect 21980 34692 22036 34702
rect 22036 34636 22148 34692
rect 21980 34560 22036 34636
rect 21756 34514 21812 34524
rect 21644 33908 21700 33918
rect 21644 32786 21700 33852
rect 21644 32734 21646 32786
rect 21698 32734 21700 32786
rect 21644 32722 21700 32734
rect 21420 32564 21476 32574
rect 21420 32470 21476 32508
rect 21756 32562 21812 32574
rect 21756 32510 21758 32562
rect 21810 32510 21812 32562
rect 20972 31714 21028 31724
rect 21756 31556 21812 32510
rect 21980 31556 22036 31566
rect 21756 31554 22036 31556
rect 21756 31502 21982 31554
rect 22034 31502 22036 31554
rect 21756 31500 22036 31502
rect 21644 30212 21700 30222
rect 21644 30118 21700 30156
rect 20860 30100 20916 30110
rect 20860 29540 20916 30044
rect 20860 29474 20916 29484
rect 21868 29876 21924 29886
rect 20524 27682 20580 27692
rect 21868 27412 21924 29820
rect 21980 27636 22036 31500
rect 22092 29988 22148 34636
rect 22316 33348 22372 33358
rect 22204 32564 22260 32574
rect 22204 32470 22260 32508
rect 22092 29764 22148 29932
rect 22316 29876 22372 33292
rect 22540 32786 22596 35196
rect 22540 32734 22542 32786
rect 22594 32734 22596 32786
rect 22540 32722 22596 32734
rect 22652 32562 22708 32574
rect 22652 32510 22654 32562
rect 22706 32510 22708 32562
rect 22652 32452 22708 32510
rect 22652 32386 22708 32396
rect 22764 30100 22820 38612
rect 23100 37828 23156 37838
rect 22876 36260 22932 36270
rect 22876 36166 22932 36204
rect 22988 35028 23044 35038
rect 22988 34934 23044 34972
rect 23100 34804 23156 37772
rect 23548 36932 23604 46396
rect 23996 45220 24052 54236
rect 24556 52834 24612 52846
rect 24556 52782 24558 52834
rect 24610 52782 24612 52834
rect 24108 52724 24164 52734
rect 24108 52630 24164 52668
rect 24556 52052 24612 52782
rect 25340 52724 25396 56028
rect 26796 56084 26852 56094
rect 26796 55990 26852 56028
rect 27804 54404 27860 54414
rect 27468 54402 27860 54404
rect 27468 54350 27806 54402
rect 27858 54350 27860 54402
rect 27468 54348 27860 54350
rect 27468 53842 27524 54348
rect 27468 53790 27470 53842
rect 27522 53790 27524 53842
rect 27468 53778 27524 53790
rect 27356 53620 27412 53630
rect 27804 53620 27860 54348
rect 27356 53526 27412 53564
rect 27692 53564 27804 53620
rect 27356 52836 27412 52846
rect 25340 52658 25396 52668
rect 25900 52724 25956 52734
rect 24556 51986 24612 51996
rect 25228 52052 25284 52062
rect 25228 50428 25284 51996
rect 25228 50372 25396 50428
rect 24556 46562 24612 46574
rect 24556 46510 24558 46562
rect 24610 46510 24612 46562
rect 24108 46450 24164 46462
rect 24108 46398 24110 46450
rect 24162 46398 24164 46450
rect 24108 46340 24164 46398
rect 24556 46452 24612 46510
rect 24556 46386 24612 46396
rect 24108 46274 24164 46284
rect 24892 45220 24948 45230
rect 23996 45164 24164 45220
rect 23884 44882 23940 44894
rect 23884 44830 23886 44882
rect 23938 44830 23940 44882
rect 23772 41746 23828 41758
rect 23772 41694 23774 41746
rect 23826 41694 23828 41746
rect 23660 40628 23716 40638
rect 23660 40534 23716 40572
rect 23772 39172 23828 41694
rect 23772 39106 23828 39116
rect 23548 36866 23604 36876
rect 23548 36370 23604 36382
rect 23548 36318 23550 36370
rect 23602 36318 23604 36370
rect 23436 36260 23492 36270
rect 22988 34748 23156 34804
rect 23324 36258 23492 36260
rect 23324 36206 23438 36258
rect 23490 36206 23492 36258
rect 23324 36204 23492 36206
rect 22876 32562 22932 32574
rect 22876 32510 22878 32562
rect 22930 32510 22932 32562
rect 22876 32340 22932 32510
rect 22876 32274 22932 32284
rect 22764 30034 22820 30044
rect 22316 29810 22372 29820
rect 22092 29698 22148 29708
rect 22204 29652 22260 29662
rect 22204 29316 22260 29596
rect 22652 29426 22708 29438
rect 22652 29374 22654 29426
rect 22706 29374 22708 29426
rect 22652 29316 22708 29374
rect 22204 29314 22708 29316
rect 22204 29262 22206 29314
rect 22258 29262 22708 29314
rect 22204 29260 22708 29262
rect 22204 29250 22260 29260
rect 21980 27570 22036 27580
rect 21868 27356 22260 27412
rect 19628 27076 19684 27086
rect 20188 27056 20244 27132
rect 21868 27188 21924 27198
rect 19628 26982 19684 27020
rect 19516 26898 19572 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 25284 19684 25294
rect 19628 24948 19684 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19740 24948 19796 24958
rect 19628 24946 19796 24948
rect 19628 24894 19742 24946
rect 19794 24894 19796 24946
rect 19628 24892 19796 24894
rect 19740 24882 19796 24892
rect 21756 24948 21812 24958
rect 21868 24948 21924 27132
rect 21756 24946 21924 24948
rect 21756 24894 21758 24946
rect 21810 24894 21924 24946
rect 21756 24892 21924 24894
rect 21756 24882 21812 24892
rect 19628 24612 19684 24622
rect 19628 24518 19684 24556
rect 21868 24612 21924 24892
rect 21868 24546 21924 24556
rect 18620 23998 18622 24050
rect 18674 23998 18676 24050
rect 18620 23492 18676 23998
rect 21196 23716 21252 23726
rect 19836 23548 20100 23558
rect 18620 23426 18676 23436
rect 19180 23492 19236 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18172 23314 18228 23324
rect 18844 23380 18900 23390
rect 18844 23286 18900 23324
rect 19180 23378 19236 23436
rect 19180 23326 19182 23378
rect 19234 23326 19236 23378
rect 19180 23314 19236 23326
rect 21196 23378 21252 23660
rect 21644 23716 21700 23726
rect 22092 23716 22148 23726
rect 21644 23622 21700 23660
rect 21980 23714 22148 23716
rect 21980 23662 22094 23714
rect 22146 23662 22148 23714
rect 21980 23660 22148 23662
rect 21196 23326 21198 23378
rect 21250 23326 21252 23378
rect 21196 23314 21252 23326
rect 17948 23214 17950 23266
rect 18002 23214 18004 23266
rect 17948 23202 18004 23214
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17836 23090 17892 23102
rect 18396 23154 18452 23166
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 16940 23044 16996 23054
rect 16940 22950 16996 22988
rect 18396 23044 18452 23102
rect 18396 22978 18452 22988
rect 21644 23044 21700 23054
rect 21644 22950 21700 22988
rect 21980 23044 22036 23660
rect 22092 23650 22148 23660
rect 22092 23380 22148 23390
rect 22204 23380 22260 27356
rect 22316 27300 22372 29260
rect 22988 28418 23044 34748
rect 23324 34690 23380 36204
rect 23436 36194 23492 36204
rect 23548 36260 23604 36318
rect 23324 34638 23326 34690
rect 23378 34638 23380 34690
rect 23324 34580 23380 34638
rect 23324 34514 23380 34524
rect 23324 32450 23380 32462
rect 23324 32398 23326 32450
rect 23378 32398 23380 32450
rect 23324 32340 23380 32398
rect 23324 32274 23380 32284
rect 23548 29540 23604 36204
rect 23660 35138 23716 35150
rect 23660 35086 23662 35138
rect 23714 35086 23716 35138
rect 23660 31890 23716 35086
rect 23772 34690 23828 34702
rect 23772 34638 23774 34690
rect 23826 34638 23828 34690
rect 23772 34244 23828 34638
rect 23772 34178 23828 34188
rect 23884 34132 23940 44830
rect 23996 43316 24052 43326
rect 23996 43222 24052 43260
rect 24108 40068 24164 45164
rect 24332 45108 24388 45118
rect 24332 44996 24388 45052
rect 24332 44994 24500 44996
rect 24332 44942 24334 44994
rect 24386 44942 24500 44994
rect 24332 44940 24500 44942
rect 24332 44930 24388 44940
rect 24332 43652 24388 43662
rect 24332 43558 24388 43596
rect 24220 41858 24276 41870
rect 24220 41806 24222 41858
rect 24274 41806 24276 41858
rect 24220 40180 24276 41806
rect 24220 40114 24276 40124
rect 24332 40964 24388 40974
rect 24108 40002 24164 40012
rect 24108 38052 24164 38062
rect 24108 37826 24164 37996
rect 24108 37774 24110 37826
rect 24162 37774 24164 37826
rect 24108 37380 24164 37774
rect 24108 37314 24164 37324
rect 24108 36372 24164 36382
rect 24108 36278 24164 36316
rect 24220 34692 24276 34702
rect 24220 34598 24276 34636
rect 23884 34066 23940 34076
rect 23996 33460 24052 33470
rect 24332 33460 24388 40908
rect 24444 38668 24500 44940
rect 24892 43764 24948 45164
rect 24892 43650 24948 43708
rect 24892 43598 24894 43650
rect 24946 43598 24948 43650
rect 24892 43586 24948 43598
rect 24668 42196 24724 42206
rect 24668 41970 24724 42140
rect 24668 41918 24670 41970
rect 24722 41918 24724 41970
rect 24668 41906 24724 41918
rect 24444 38612 24948 38668
rect 24556 38164 24612 38174
rect 24556 38070 24612 38108
rect 24444 36932 24500 36942
rect 24444 33684 24500 36876
rect 24892 36594 24948 38612
rect 25004 37828 25060 37838
rect 25004 37734 25060 37772
rect 25004 37380 25060 37390
rect 25004 37286 25060 37324
rect 24892 36542 24894 36594
rect 24946 36542 24948 36594
rect 24892 36530 24948 36542
rect 25116 36484 25172 36494
rect 24892 36372 24948 36382
rect 24780 36260 24836 36270
rect 24780 36166 24836 36204
rect 24892 35476 24948 36316
rect 24556 35140 24612 35150
rect 24780 35140 24836 35150
rect 24556 35138 24836 35140
rect 24556 35086 24558 35138
rect 24610 35086 24782 35138
rect 24834 35086 24836 35138
rect 24556 35084 24836 35086
rect 24556 35074 24612 35084
rect 24780 35074 24836 35084
rect 24892 34916 24948 35420
rect 25004 36258 25060 36270
rect 25004 36206 25006 36258
rect 25058 36206 25060 36258
rect 25004 35140 25060 36206
rect 25004 35074 25060 35084
rect 24668 34860 24948 34916
rect 25004 34916 25060 34926
rect 25116 34916 25172 36428
rect 25228 36482 25284 36494
rect 25228 36430 25230 36482
rect 25282 36430 25284 36482
rect 25228 36372 25284 36430
rect 25228 36306 25284 36316
rect 25340 35028 25396 50372
rect 25900 40626 25956 52668
rect 27244 52722 27300 52734
rect 27244 52670 27246 52722
rect 27298 52670 27300 52722
rect 27244 50932 27300 52670
rect 27244 50866 27300 50876
rect 27356 52164 27412 52780
rect 27580 52164 27636 52174
rect 27356 52162 27636 52164
rect 27356 52110 27582 52162
rect 27634 52110 27636 52162
rect 27356 52108 27636 52110
rect 26572 48244 26628 48254
rect 26348 40740 26404 40750
rect 26348 40628 26404 40684
rect 25900 40574 25902 40626
rect 25954 40574 25956 40626
rect 25900 40516 25956 40574
rect 25900 40450 25956 40460
rect 26236 40626 26404 40628
rect 26236 40574 26350 40626
rect 26402 40574 26404 40626
rect 26236 40572 26404 40574
rect 26012 39396 26068 39406
rect 25676 38164 25732 38174
rect 25564 38052 25620 38062
rect 25564 37958 25620 37996
rect 25676 37938 25732 38108
rect 25676 37886 25678 37938
rect 25730 37886 25732 37938
rect 25676 37874 25732 37886
rect 25900 37940 25956 37950
rect 25900 37846 25956 37884
rect 25788 37380 25844 37390
rect 26012 37380 26068 39340
rect 26124 38052 26180 38062
rect 26124 37828 26180 37996
rect 26124 37762 26180 37772
rect 25844 37324 26068 37380
rect 25676 37268 25732 37278
rect 25788 37248 25844 37324
rect 26236 37268 26292 40572
rect 26348 40562 26404 40572
rect 26348 39396 26404 39406
rect 26348 39302 26404 39340
rect 25676 37044 25732 37212
rect 25676 36978 25732 36988
rect 26012 37212 26292 37268
rect 26460 38500 26516 38510
rect 25452 36482 25508 36494
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 25452 35364 25508 36430
rect 25676 36482 25732 36494
rect 25676 36430 25678 36482
rect 25730 36430 25732 36482
rect 25676 36036 25732 36430
rect 25676 35970 25732 35980
rect 25452 35298 25508 35308
rect 26012 35588 26068 37212
rect 26236 36258 26292 36270
rect 26236 36206 26238 36258
rect 26290 36206 26292 36258
rect 26236 36036 26292 36206
rect 26236 35970 26292 35980
rect 25452 35028 25508 35038
rect 25340 35026 25508 35028
rect 25340 34974 25454 35026
rect 25506 34974 25508 35026
rect 25340 34972 25508 34974
rect 25452 34962 25508 34972
rect 25228 34916 25284 34926
rect 25116 34914 25284 34916
rect 25116 34862 25230 34914
rect 25282 34862 25284 34914
rect 25116 34860 25284 34862
rect 24444 33628 24612 33684
rect 24444 33460 24500 33470
rect 24332 33458 24500 33460
rect 24332 33406 24446 33458
rect 24498 33406 24500 33458
rect 24332 33404 24500 33406
rect 23996 33366 24052 33404
rect 24444 33348 24500 33404
rect 24444 33282 24500 33292
rect 23772 32452 23828 32462
rect 23772 32358 23828 32396
rect 23660 31838 23662 31890
rect 23714 31838 23716 31890
rect 23660 31826 23716 31838
rect 24108 32340 24164 32350
rect 23884 31666 23940 31678
rect 23884 31614 23886 31666
rect 23938 31614 23940 31666
rect 23660 31554 23716 31566
rect 23660 31502 23662 31554
rect 23714 31502 23716 31554
rect 23660 31220 23716 31502
rect 23884 31556 23940 31614
rect 23884 31490 23940 31500
rect 23660 31154 23716 31164
rect 23548 29474 23604 29484
rect 23100 29426 23156 29438
rect 23100 29374 23102 29426
rect 23154 29374 23156 29426
rect 23100 29092 23156 29374
rect 23324 29426 23380 29438
rect 23324 29374 23326 29426
rect 23378 29374 23380 29426
rect 23100 29026 23156 29036
rect 23212 29314 23268 29326
rect 23212 29262 23214 29314
rect 23266 29262 23268 29314
rect 23100 28644 23156 28654
rect 23100 28550 23156 28588
rect 22988 28366 22990 28418
rect 23042 28366 23044 28418
rect 22988 28354 23044 28366
rect 22316 24946 22372 27244
rect 22428 28084 22484 28094
rect 22428 27188 22484 28028
rect 23212 27970 23268 29262
rect 23324 29316 23380 29374
rect 23772 29316 23828 29326
rect 23324 29314 23828 29316
rect 23324 29262 23774 29314
rect 23826 29262 23828 29314
rect 23324 29260 23828 29262
rect 23436 29092 23492 29102
rect 23324 28868 23380 28878
rect 23324 28082 23380 28812
rect 23436 28644 23492 29036
rect 23436 28550 23492 28588
rect 23548 28754 23604 29260
rect 23772 29250 23828 29260
rect 23548 28702 23550 28754
rect 23602 28702 23604 28754
rect 23548 28532 23604 28702
rect 23548 28466 23604 28476
rect 23324 28030 23326 28082
rect 23378 28030 23380 28082
rect 23324 28018 23380 28030
rect 23772 27972 23828 27982
rect 23212 27918 23214 27970
rect 23266 27918 23268 27970
rect 23212 27906 23268 27918
rect 23660 27916 23772 27972
rect 23548 27858 23604 27870
rect 23548 27806 23550 27858
rect 23602 27806 23604 27858
rect 23548 27636 23604 27806
rect 23548 27570 23604 27580
rect 22428 27122 22484 27132
rect 23324 27524 23380 27534
rect 22876 27074 22932 27086
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22540 26964 22596 26974
rect 22540 25730 22596 26908
rect 22540 25678 22542 25730
rect 22594 25678 22596 25730
rect 22540 25666 22596 25678
rect 22316 24894 22318 24946
rect 22370 24894 22372 24946
rect 22316 24882 22372 24894
rect 22428 25620 22484 25630
rect 22428 24836 22484 25564
rect 22876 25284 22932 27022
rect 23212 27076 23268 27086
rect 23212 26850 23268 27020
rect 23324 27074 23380 27468
rect 23324 27022 23326 27074
rect 23378 27022 23380 27074
rect 23324 27010 23380 27022
rect 23436 27412 23492 27422
rect 23212 26798 23214 26850
rect 23266 26798 23268 26850
rect 23212 26786 23268 26798
rect 23436 26852 23492 27356
rect 23548 27076 23604 27086
rect 23660 27076 23716 27916
rect 23772 27878 23828 27916
rect 24108 27972 24164 32284
rect 24332 31556 24388 31566
rect 24332 31462 24388 31500
rect 24220 29314 24276 29326
rect 24220 29262 24222 29314
rect 24274 29262 24276 29314
rect 24220 28868 24276 29262
rect 24220 28802 24276 28812
rect 24220 28642 24276 28654
rect 24220 28590 24222 28642
rect 24274 28590 24276 28642
rect 24220 28532 24276 28590
rect 24220 28466 24276 28476
rect 24220 27972 24276 27982
rect 24164 27970 24276 27972
rect 24164 27918 24222 27970
rect 24274 27918 24276 27970
rect 24164 27916 24276 27918
rect 24108 27840 24164 27916
rect 24220 27906 24276 27916
rect 23548 27074 23716 27076
rect 23548 27022 23550 27074
rect 23602 27022 23716 27074
rect 23548 27020 23716 27022
rect 23548 27010 23604 27020
rect 23436 26796 23604 26852
rect 22988 25620 23044 25630
rect 22988 25526 23044 25564
rect 22876 25218 22932 25228
rect 23548 25060 23604 26796
rect 23660 26514 23716 27020
rect 23660 26462 23662 26514
rect 23714 26462 23716 26514
rect 23660 26450 23716 26462
rect 23996 27524 24052 27534
rect 23996 26514 24052 27468
rect 24444 27188 24500 27198
rect 24444 27074 24500 27132
rect 24556 27186 24612 33628
rect 24668 30996 24724 34860
rect 25004 34822 25060 34860
rect 25228 34692 25284 34860
rect 25452 34804 25508 34814
rect 25452 34710 25508 34748
rect 25116 34132 25172 34142
rect 25004 33124 25060 33134
rect 25004 33030 25060 33068
rect 25004 32564 25060 32574
rect 24892 32452 24948 32462
rect 25004 32452 25060 32508
rect 24892 32450 25060 32452
rect 24892 32398 24894 32450
rect 24946 32398 25060 32450
rect 24892 32396 25060 32398
rect 24892 32386 24948 32396
rect 24780 31554 24836 31566
rect 24780 31502 24782 31554
rect 24834 31502 24836 31554
rect 24780 31220 24836 31502
rect 24780 31154 24836 31164
rect 24668 30940 24836 30996
rect 24668 28644 24724 28654
rect 24668 28550 24724 28588
rect 24668 27746 24724 27758
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24668 27636 24724 27694
rect 24668 27570 24724 27580
rect 24556 27134 24558 27186
rect 24610 27134 24612 27186
rect 24556 27122 24612 27134
rect 24444 27022 24446 27074
rect 24498 27022 24500 27074
rect 24444 27010 24500 27022
rect 24780 27074 24836 30940
rect 24892 29652 24948 29662
rect 24892 29558 24948 29596
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24668 26964 24724 27002
rect 24668 26898 24724 26908
rect 23996 26462 23998 26514
rect 24050 26462 24052 26514
rect 23996 25732 24052 26462
rect 24556 26516 24612 26526
rect 24780 26516 24836 27022
rect 25004 26908 25060 32396
rect 25116 27412 25172 34076
rect 25228 33684 25284 34636
rect 25228 33618 25284 33628
rect 25676 34690 25732 34702
rect 25676 34638 25678 34690
rect 25730 34638 25732 34690
rect 25676 34244 25732 34638
rect 25452 33460 25508 33470
rect 25452 33366 25508 33404
rect 25564 33234 25620 33246
rect 25564 33182 25566 33234
rect 25618 33182 25620 33234
rect 25564 33124 25620 33182
rect 25564 33058 25620 33068
rect 25676 32676 25732 34188
rect 26012 33460 26068 35532
rect 26236 35364 26292 35374
rect 26012 33394 26068 33404
rect 26124 34020 26180 34030
rect 25788 33348 25844 33358
rect 25788 33254 25844 33292
rect 26124 33346 26180 33964
rect 26124 33294 26126 33346
rect 26178 33294 26180 33346
rect 25676 32610 25732 32620
rect 26012 32562 26068 32574
rect 26012 32510 26014 32562
rect 26066 32510 26068 32562
rect 26012 32340 26068 32510
rect 26012 32274 26068 32284
rect 25340 30884 25396 30894
rect 25116 27346 25172 27356
rect 25228 28644 25284 28654
rect 25116 27076 25172 27086
rect 25116 26982 25172 27020
rect 24556 26514 24836 26516
rect 24556 26462 24558 26514
rect 24610 26462 24836 26514
rect 24556 26460 24836 26462
rect 24892 26852 25060 26908
rect 25228 26964 25284 28588
rect 25340 27298 25396 30828
rect 26124 30212 26180 33294
rect 26236 32788 26292 35308
rect 26348 34916 26404 34926
rect 26348 34244 26404 34860
rect 26348 34178 26404 34188
rect 26460 33570 26516 38444
rect 26572 38274 26628 48188
rect 26796 47572 26852 47582
rect 26796 47478 26852 47516
rect 27356 47572 27412 52108
rect 27580 52098 27636 52108
rect 27692 49250 27748 53564
rect 27804 53554 27860 53564
rect 28252 53508 28308 53518
rect 28140 53506 28308 53508
rect 28140 53454 28254 53506
rect 28306 53454 28308 53506
rect 28140 53452 28308 53454
rect 28028 53060 28084 53070
rect 28140 53060 28196 53452
rect 28252 53442 28308 53452
rect 28084 53004 28196 53060
rect 28252 53060 28308 53070
rect 28364 53060 28420 56140
rect 29260 56082 29316 56094
rect 29260 56030 29262 56082
rect 29314 56030 29316 56082
rect 28588 55970 28644 55982
rect 28588 55918 28590 55970
rect 28642 55918 28644 55970
rect 28588 55188 28644 55918
rect 28588 55122 28644 55132
rect 29260 55188 29316 56030
rect 29932 55970 29988 56590
rect 31388 56308 31444 56318
rect 31500 56308 31556 59200
rect 31388 56306 31556 56308
rect 31388 56254 31390 56306
rect 31442 56254 31556 56306
rect 31388 56252 31556 56254
rect 31388 56242 31444 56252
rect 31500 56084 31556 56252
rect 34748 56308 34804 56318
rect 34860 56308 34916 59200
rect 37436 56308 37492 56318
rect 37548 56308 37604 59200
rect 34748 56306 35252 56308
rect 34748 56254 34750 56306
rect 34802 56254 35252 56306
rect 34748 56252 35252 56254
rect 34748 56242 34804 56252
rect 31836 56196 31892 56206
rect 31836 56102 31892 56140
rect 35196 56194 35252 56252
rect 37436 56306 37940 56308
rect 37436 56254 37438 56306
rect 37490 56254 37940 56306
rect 37436 56252 37940 56254
rect 37436 56242 37492 56252
rect 35196 56142 35198 56194
rect 35250 56142 35252 56194
rect 35196 56130 35252 56142
rect 35532 56194 35588 56206
rect 35532 56142 35534 56194
rect 35586 56142 35588 56194
rect 31500 56018 31556 56028
rect 32060 56084 32116 56094
rect 32060 55990 32116 56028
rect 29932 55918 29934 55970
rect 29986 55918 29988 55970
rect 29932 55906 29988 55918
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35532 55468 35588 56142
rect 37884 56194 37940 56252
rect 37884 56142 37886 56194
rect 37938 56142 37940 56194
rect 37884 56130 37940 56142
rect 38220 56196 38276 56206
rect 38220 56102 38276 56140
rect 39788 56196 39844 56206
rect 35532 55412 35812 55468
rect 29260 55122 29316 55132
rect 28252 53058 28420 53060
rect 28252 53006 28254 53058
rect 28306 53006 28420 53058
rect 28252 53004 28420 53006
rect 28476 54628 28532 54638
rect 28028 52966 28084 53004
rect 28252 52994 28308 53004
rect 27916 52724 27972 52734
rect 27692 49198 27694 49250
rect 27746 49198 27748 49250
rect 27692 48354 27748 49198
rect 27692 48302 27694 48354
rect 27746 48302 27748 48354
rect 27692 48290 27748 48302
rect 27804 52722 27972 52724
rect 27804 52670 27918 52722
rect 27970 52670 27972 52722
rect 27804 52668 27972 52670
rect 27580 48020 27636 48030
rect 27356 47478 27412 47516
rect 27468 48018 27636 48020
rect 27468 47966 27582 48018
rect 27634 47966 27636 48018
rect 27468 47964 27636 47966
rect 27244 47234 27300 47246
rect 27244 47182 27246 47234
rect 27298 47182 27300 47234
rect 27244 42196 27300 47182
rect 27468 43708 27524 47964
rect 27580 47954 27636 47964
rect 27804 47572 27860 52668
rect 27916 52658 27972 52668
rect 28476 52500 28532 54572
rect 29148 54402 29204 54414
rect 29148 54350 29150 54402
rect 29202 54350 29204 54402
rect 28700 54292 28756 54302
rect 28700 53730 28756 54236
rect 28700 53678 28702 53730
rect 28754 53678 28756 53730
rect 28700 53666 28756 53678
rect 28812 53620 28868 53630
rect 28812 53526 28868 53564
rect 29148 53620 29204 54350
rect 30716 54402 30772 54414
rect 30716 54350 30718 54402
rect 30770 54350 30772 54402
rect 30268 53956 30324 53966
rect 30268 53862 30324 53900
rect 29148 53554 29204 53564
rect 29484 53620 29540 53630
rect 29484 53506 29540 53564
rect 30380 53620 30436 53630
rect 30380 53526 30436 53564
rect 30716 53620 30772 54350
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 32508 53732 32564 53742
rect 32508 53638 32564 53676
rect 32620 53732 32676 53742
rect 33068 53732 33124 53742
rect 32620 53730 33124 53732
rect 32620 53678 32622 53730
rect 32674 53678 33070 53730
rect 33122 53678 33124 53730
rect 32620 53676 33124 53678
rect 30716 53554 30772 53564
rect 31052 53620 31108 53630
rect 29484 53454 29486 53506
rect 29538 53454 29540 53506
rect 29036 53172 29092 53182
rect 29036 53078 29092 53116
rect 28252 52444 28532 52500
rect 29148 52834 29204 52846
rect 29148 52782 29150 52834
rect 29202 52782 29204 52834
rect 27580 47516 27860 47572
rect 27916 49250 27972 49262
rect 27916 49198 27918 49250
rect 27970 49198 27972 49250
rect 27916 49138 27972 49198
rect 27916 49086 27918 49138
rect 27970 49086 27972 49138
rect 27580 45332 27636 47516
rect 27916 47460 27972 49086
rect 28028 47460 28084 47470
rect 27916 47458 28084 47460
rect 27916 47406 28030 47458
rect 28082 47406 28084 47458
rect 27916 47404 28084 47406
rect 27916 47236 27972 47246
rect 27916 47142 27972 47180
rect 28028 47012 28084 47404
rect 28252 47348 28308 52444
rect 28476 52276 28532 52286
rect 28476 52182 28532 52220
rect 29148 52276 29204 52782
rect 29148 52210 29204 52220
rect 29484 52276 29540 53454
rect 30492 53508 30548 53518
rect 29708 53284 29764 53294
rect 29708 53170 29764 53228
rect 29708 53118 29710 53170
rect 29762 53118 29764 53170
rect 29708 53106 29764 53118
rect 30492 53060 30548 53452
rect 30940 53506 30996 53518
rect 30940 53454 30942 53506
rect 30994 53454 30996 53506
rect 30492 53058 30772 53060
rect 30492 53006 30494 53058
rect 30546 53006 30772 53058
rect 30492 53004 30772 53006
rect 30492 52994 30548 53004
rect 29820 52836 29876 52846
rect 29820 52276 29876 52780
rect 30380 52722 30436 52734
rect 30380 52670 30382 52722
rect 30434 52670 30436 52722
rect 30044 52276 30100 52286
rect 29820 52220 30044 52276
rect 29484 52182 29540 52220
rect 28364 52164 28420 52174
rect 30044 52144 30100 52220
rect 28364 52070 28420 52108
rect 30380 51380 30436 52670
rect 30716 52274 30772 53004
rect 30940 52948 30996 53454
rect 31052 53060 31108 53564
rect 31500 53506 31556 53518
rect 31500 53454 31502 53506
rect 31554 53454 31556 53506
rect 31164 53060 31220 53070
rect 31500 53060 31556 53454
rect 31052 53058 31556 53060
rect 31052 53006 31166 53058
rect 31218 53006 31556 53058
rect 31052 53004 31556 53006
rect 31164 52994 31220 53004
rect 30940 52882 30996 52892
rect 31500 52948 31556 53004
rect 31612 52948 31668 52958
rect 31500 52946 31668 52948
rect 31500 52894 31614 52946
rect 31666 52894 31668 52946
rect 31500 52892 31668 52894
rect 30716 52222 30718 52274
rect 30770 52222 30772 52274
rect 30716 52164 30772 52222
rect 30716 52098 30772 52108
rect 31052 52722 31108 52734
rect 31052 52670 31054 52722
rect 31106 52670 31108 52722
rect 31052 51492 31108 52670
rect 31388 52612 31444 52622
rect 31388 52386 31444 52556
rect 31388 52334 31390 52386
rect 31442 52334 31444 52386
rect 31388 52322 31444 52334
rect 31500 52274 31556 52892
rect 31612 52882 31668 52892
rect 32620 52276 32676 53676
rect 33068 53666 33124 53676
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 31500 52222 31502 52274
rect 31554 52222 31556 52274
rect 31500 52164 31556 52222
rect 32508 52220 32620 52276
rect 31500 52108 32004 52164
rect 31052 51426 31108 51436
rect 31948 51938 32004 52108
rect 31948 51886 31950 51938
rect 32002 51886 32004 51938
rect 30380 51314 30436 51324
rect 29820 51156 29876 51166
rect 27804 46956 28028 47012
rect 27804 46786 27860 46956
rect 28028 46946 28084 46956
rect 28140 47292 28308 47348
rect 28364 49700 28420 49710
rect 27804 46734 27806 46786
rect 27858 46734 27860 46786
rect 27804 46722 27860 46734
rect 27580 45200 27636 45276
rect 27692 46450 27748 46462
rect 27692 46398 27694 46450
rect 27746 46398 27748 46450
rect 27468 43652 27636 43708
rect 27244 42130 27300 42140
rect 26796 41076 26852 41086
rect 26796 40628 26852 41020
rect 26572 38222 26574 38274
rect 26626 38222 26628 38274
rect 26572 38210 26628 38222
rect 26684 40626 26852 40628
rect 26684 40574 26798 40626
rect 26850 40574 26852 40626
rect 26684 40572 26852 40574
rect 26684 38052 26740 40572
rect 26796 40562 26852 40572
rect 27244 40516 27300 40526
rect 26908 40292 26964 40302
rect 26908 39732 26964 40236
rect 27244 39732 27300 40460
rect 27468 40516 27524 40526
rect 27468 40422 27524 40460
rect 27356 40292 27412 40302
rect 27356 40198 27412 40236
rect 27580 39844 27636 43652
rect 27692 40628 27748 46398
rect 27916 44996 27972 45006
rect 27916 44902 27972 44940
rect 27916 41076 27972 41086
rect 27692 40562 27748 40572
rect 27804 40740 27860 40750
rect 27804 40514 27860 40684
rect 27804 40462 27806 40514
rect 27858 40462 27860 40514
rect 27804 40450 27860 40462
rect 27916 40628 27972 41020
rect 27916 40402 27972 40572
rect 27916 40350 27918 40402
rect 27970 40350 27972 40402
rect 27916 40338 27972 40350
rect 28140 40292 28196 47292
rect 28252 47012 28308 47022
rect 28252 46898 28308 46956
rect 28252 46846 28254 46898
rect 28306 46846 28308 46898
rect 28252 46834 28308 46846
rect 28364 43708 28420 49644
rect 29596 48804 29652 48814
rect 28700 48132 28756 48142
rect 29148 48132 29204 48142
rect 28700 48130 29204 48132
rect 28700 48078 28702 48130
rect 28754 48078 29150 48130
rect 29202 48078 29204 48130
rect 28700 48076 29204 48078
rect 28700 48066 28756 48076
rect 28588 48018 28644 48030
rect 28588 47966 28590 48018
rect 28642 47966 28644 48018
rect 28588 47684 28644 47966
rect 28476 47628 28644 47684
rect 28476 46900 28532 47628
rect 28700 47348 28756 47358
rect 28924 47348 28980 48076
rect 29148 48066 29204 48076
rect 28700 47346 28980 47348
rect 28700 47294 28702 47346
rect 28754 47294 28980 47346
rect 28700 47292 28980 47294
rect 28588 47234 28644 47246
rect 28588 47182 28590 47234
rect 28642 47182 28644 47234
rect 28588 47124 28644 47182
rect 28588 47058 28644 47068
rect 28700 47012 28756 47292
rect 28476 46844 28644 46900
rect 28588 45220 28644 46844
rect 28700 46898 28756 46956
rect 28700 46846 28702 46898
rect 28754 46846 28756 46898
rect 28700 46834 28756 46846
rect 29484 47234 29540 47246
rect 29484 47182 29486 47234
rect 29538 47182 29540 47234
rect 29484 47012 29540 47182
rect 29484 46786 29540 46956
rect 29484 46734 29486 46786
rect 29538 46734 29540 46786
rect 29484 46722 29540 46734
rect 29372 46564 29428 46574
rect 29372 46470 29428 46508
rect 28588 45154 28644 45164
rect 28700 45666 28756 45678
rect 28700 45614 28702 45666
rect 28754 45614 28756 45666
rect 28700 45108 28756 45614
rect 28700 45042 28756 45052
rect 29260 45332 29316 45342
rect 29260 45106 29316 45276
rect 29260 45054 29262 45106
rect 29314 45054 29316 45106
rect 29260 45042 29316 45054
rect 28588 44994 28644 45006
rect 28588 44942 28590 44994
rect 28642 44942 28644 44994
rect 28140 40226 28196 40236
rect 28252 43652 28420 43708
rect 28476 44882 28532 44894
rect 28476 44830 28478 44882
rect 28530 44830 28532 44882
rect 26796 39676 26964 39732
rect 27020 39730 27300 39732
rect 27020 39678 27246 39730
rect 27298 39678 27300 39730
rect 27020 39676 27300 39678
rect 26796 39396 26852 39676
rect 26796 39302 26852 39340
rect 27020 39060 27076 39676
rect 27244 39666 27300 39676
rect 27356 39788 27636 39844
rect 27356 39620 27412 39788
rect 28252 39732 28308 43652
rect 28476 42644 28532 44830
rect 28588 44436 28644 44942
rect 29484 44882 29540 44894
rect 29484 44830 29486 44882
rect 29538 44830 29540 44882
rect 28812 44436 28868 44446
rect 28588 44380 28812 44436
rect 28812 44342 28868 44380
rect 28476 42578 28532 42588
rect 29484 42196 29540 44830
rect 29596 44548 29652 48748
rect 29596 44482 29652 44492
rect 29708 45108 29764 45118
rect 29484 42130 29540 42140
rect 28364 41300 28420 41310
rect 28364 40626 28420 41244
rect 28812 41300 28868 41310
rect 28812 41206 28868 41244
rect 29708 41188 29764 45052
rect 29708 41122 29764 41132
rect 29820 41300 29876 51100
rect 30380 49924 30436 49934
rect 31948 49924 32004 51886
rect 32396 50370 32452 50382
rect 32396 50318 32398 50370
rect 32450 50318 32452 50370
rect 32172 49924 32228 49934
rect 31948 49868 32172 49924
rect 29932 47012 29988 47022
rect 29932 46898 29988 46956
rect 29932 46846 29934 46898
rect 29986 46846 29988 46898
rect 29932 46834 29988 46846
rect 29932 45332 29988 45342
rect 29932 45238 29988 45276
rect 30268 45220 30324 45230
rect 30156 45106 30212 45118
rect 30156 45054 30158 45106
rect 30210 45054 30212 45106
rect 29932 44996 29988 45006
rect 29932 41300 29988 44940
rect 30044 44994 30100 45006
rect 30044 44942 30046 44994
rect 30098 44942 30100 44994
rect 30044 43652 30100 44942
rect 30156 44996 30212 45054
rect 30156 44930 30212 44940
rect 30156 44548 30212 44558
rect 30156 44454 30212 44492
rect 30268 44436 30324 45164
rect 30380 45108 30436 49868
rect 31500 49700 31556 49710
rect 31388 49586 31444 49598
rect 31388 49534 31390 49586
rect 31442 49534 31444 49586
rect 31388 48468 31444 49534
rect 31388 48402 31444 48412
rect 31500 46004 31556 49644
rect 32172 49700 32228 49868
rect 32396 49924 32452 50318
rect 32396 49858 32452 49868
rect 32172 49634 32228 49644
rect 32060 49588 32116 49598
rect 32060 49494 32116 49532
rect 31948 49140 32004 49150
rect 32396 49140 32452 49150
rect 32508 49140 32564 52220
rect 32620 52210 32676 52220
rect 35532 52164 35588 52174
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35532 50706 35588 52108
rect 35532 50654 35534 50706
rect 35586 50654 35588 50706
rect 35532 50642 35588 50654
rect 32620 49924 32676 49934
rect 32620 49830 32676 49868
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 31948 49138 32508 49140
rect 31948 49086 31950 49138
rect 32002 49086 32398 49138
rect 32450 49086 32508 49138
rect 31948 49084 32508 49086
rect 31948 49074 32004 49084
rect 31836 48916 31892 48926
rect 31836 48822 31892 48860
rect 31276 45948 31556 46004
rect 31612 47460 31668 47470
rect 30716 45892 30772 45902
rect 30716 45798 30772 45836
rect 31164 45892 31220 45902
rect 30604 45668 30660 45678
rect 30380 45042 30436 45052
rect 30492 45666 30660 45668
rect 30492 45614 30606 45666
rect 30658 45614 30660 45666
rect 30492 45612 30660 45614
rect 30268 44304 30324 44380
rect 30044 43586 30100 43596
rect 30492 42980 30548 45612
rect 30604 45602 30660 45612
rect 31164 45666 31220 45836
rect 31164 45614 31166 45666
rect 31218 45614 31220 45666
rect 30940 45444 30996 45454
rect 30716 45332 30772 45342
rect 30716 45238 30772 45276
rect 30604 45220 30660 45230
rect 30604 43762 30660 45164
rect 30604 43710 30606 43762
rect 30658 43710 30660 43762
rect 30604 43698 30660 43710
rect 30828 45108 30884 45118
rect 30828 43708 30884 45052
rect 30492 42914 30548 42924
rect 30716 43652 30884 43708
rect 30156 41300 30212 41310
rect 29932 41244 30156 41300
rect 29596 41076 29652 41086
rect 28364 40574 28366 40626
rect 28418 40574 28420 40626
rect 28364 40562 28420 40574
rect 28924 41074 29652 41076
rect 28924 41022 29598 41074
rect 29650 41022 29652 41074
rect 28924 41020 29652 41022
rect 28476 40516 28532 40526
rect 27356 39554 27412 39564
rect 27468 39676 28308 39732
rect 28364 40292 28420 40302
rect 27020 38946 27076 39004
rect 27020 38894 27022 38946
rect 27074 38894 27076 38946
rect 27020 38882 27076 38894
rect 26684 37986 26740 37996
rect 26908 38610 26964 38622
rect 26908 38558 26910 38610
rect 26962 38558 26964 38610
rect 26908 37828 26964 38558
rect 26684 37826 26964 37828
rect 26684 37774 26910 37826
rect 26962 37774 26964 37826
rect 26684 37772 26964 37774
rect 26572 37154 26628 37166
rect 26572 37102 26574 37154
rect 26626 37102 26628 37154
rect 26572 37044 26628 37102
rect 26572 36978 26628 36988
rect 26572 36260 26628 36270
rect 26572 34244 26628 36204
rect 26684 35026 26740 37772
rect 26908 37268 26964 37772
rect 27356 38276 27412 38286
rect 27356 37940 27412 38220
rect 27356 37826 27412 37884
rect 27356 37774 27358 37826
rect 27410 37774 27412 37826
rect 27356 37490 27412 37774
rect 27356 37438 27358 37490
rect 27410 37438 27412 37490
rect 27356 37426 27412 37438
rect 26908 37202 26964 37212
rect 27244 37380 27300 37390
rect 27132 36596 27188 36606
rect 27244 36596 27300 37324
rect 27132 36594 27300 36596
rect 27132 36542 27134 36594
rect 27186 36542 27300 36594
rect 27132 36540 27300 36542
rect 27132 36530 27188 36540
rect 26684 34974 26686 35026
rect 26738 34974 26740 35026
rect 26684 34804 26740 34974
rect 26684 34738 26740 34748
rect 26908 35140 26964 35150
rect 26572 34188 26740 34244
rect 26572 34020 26628 34030
rect 26572 33926 26628 33964
rect 26460 33518 26462 33570
rect 26514 33518 26516 33570
rect 26460 33506 26516 33518
rect 26684 33348 26740 34188
rect 26460 33292 26740 33348
rect 26348 32788 26404 32798
rect 26236 32786 26404 32788
rect 26236 32734 26350 32786
rect 26402 32734 26404 32786
rect 26236 32732 26404 32734
rect 26348 32722 26404 32732
rect 26236 32564 26292 32574
rect 26236 32470 26292 32508
rect 26124 30146 26180 30156
rect 25676 29652 25732 29662
rect 25676 29558 25732 29596
rect 26236 29540 26292 29550
rect 26460 29540 26516 33292
rect 26796 33236 26852 33246
rect 26684 33234 26852 33236
rect 26684 33182 26798 33234
rect 26850 33182 26852 33234
rect 26684 33180 26852 33182
rect 26908 33236 26964 35084
rect 27020 34020 27076 34030
rect 27020 34018 27188 34020
rect 27020 33966 27022 34018
rect 27074 33966 27188 34018
rect 27020 33964 27188 33966
rect 27020 33954 27076 33964
rect 27020 33236 27076 33246
rect 26908 33234 27076 33236
rect 26908 33182 27022 33234
rect 27074 33182 27076 33234
rect 26908 33180 27076 33182
rect 26684 32562 26740 33180
rect 26796 33170 26852 33180
rect 27020 33170 27076 33180
rect 27132 33234 27188 33964
rect 27468 33236 27524 39676
rect 28364 39618 28420 40236
rect 28364 39566 28366 39618
rect 28418 39566 28420 39618
rect 28364 39554 28420 39566
rect 28476 39618 28532 40460
rect 28700 39732 28756 39742
rect 28924 39732 28980 41020
rect 29596 41010 29652 41020
rect 29820 41074 29876 41244
rect 29820 41022 29822 41074
rect 29874 41022 29876 41074
rect 29820 41010 29876 41022
rect 29932 41076 29988 41086
rect 29708 40962 29764 40974
rect 29708 40910 29710 40962
rect 29762 40910 29764 40962
rect 29708 40292 29764 40910
rect 29708 40226 29764 40236
rect 28700 39730 28980 39732
rect 28700 39678 28702 39730
rect 28754 39678 28980 39730
rect 28700 39676 28980 39678
rect 28700 39666 28756 39676
rect 28476 39566 28478 39618
rect 28530 39566 28532 39618
rect 28476 39554 28532 39566
rect 28812 39506 28868 39518
rect 28812 39454 28814 39506
rect 28866 39454 28868 39506
rect 27804 39394 27860 39406
rect 27804 39342 27806 39394
rect 27858 39342 27860 39394
rect 27580 39060 27636 39070
rect 27580 38966 27636 39004
rect 27804 38388 27860 39342
rect 27804 38322 27860 38332
rect 28812 38388 28868 39454
rect 28812 38322 28868 38332
rect 28812 37268 28868 37278
rect 28812 37174 28868 37212
rect 29148 37266 29204 37278
rect 29148 37214 29150 37266
rect 29202 37214 29204 37266
rect 29148 37044 29204 37214
rect 29148 36978 29204 36988
rect 29708 36260 29764 36270
rect 29708 36166 29764 36204
rect 29708 35812 29764 35822
rect 29708 35718 29764 35756
rect 29932 35812 29988 41020
rect 30044 40628 30100 40638
rect 30044 40534 30100 40572
rect 30156 40404 30212 41244
rect 30044 40348 30212 40404
rect 30492 40516 30548 40526
rect 30492 40402 30548 40460
rect 30492 40350 30494 40402
rect 30546 40350 30548 40402
rect 30044 36260 30100 40348
rect 30044 36194 30100 36204
rect 30156 39060 30212 39070
rect 30156 37938 30212 39004
rect 30492 38276 30548 40350
rect 30716 38668 30772 43652
rect 30940 39396 30996 45388
rect 31164 45220 31220 45614
rect 31164 45154 31220 45164
rect 31164 44436 31220 44446
rect 31276 44436 31332 45948
rect 31500 45444 31556 45454
rect 31500 45218 31556 45388
rect 31500 45166 31502 45218
rect 31554 45166 31556 45218
rect 31500 45154 31556 45166
rect 31388 44884 31444 44894
rect 31388 44790 31444 44828
rect 31164 44434 31332 44436
rect 31164 44382 31166 44434
rect 31218 44382 31332 44434
rect 31164 44380 31332 44382
rect 31164 44370 31220 44380
rect 31052 44324 31108 44334
rect 31052 44230 31108 44268
rect 31276 43652 31332 44380
rect 31612 44436 31668 47404
rect 31724 47012 31780 47022
rect 31724 46002 31780 46956
rect 31724 45950 31726 46002
rect 31778 45950 31780 46002
rect 31724 45444 31780 45950
rect 32396 46004 32452 49084
rect 32508 49008 32564 49084
rect 35756 48916 35812 55412
rect 38444 54740 38500 54750
rect 35980 54404 36036 54414
rect 35868 49924 35924 49934
rect 35868 49830 35924 49868
rect 35980 49700 36036 54348
rect 38444 53956 38500 54684
rect 38892 53956 38948 53966
rect 38444 53954 38948 53956
rect 38444 53902 38894 53954
rect 38946 53902 38948 53954
rect 38444 53900 38948 53902
rect 38444 53730 38500 53900
rect 38892 53890 38948 53900
rect 39788 53954 39844 56140
rect 41132 56196 41188 59200
rect 46284 56420 46340 59200
rect 46284 56364 46900 56420
rect 46172 56308 46228 56318
rect 46284 56308 46340 56364
rect 46172 56306 46340 56308
rect 46172 56254 46174 56306
rect 46226 56254 46340 56306
rect 46172 56252 46340 56254
rect 46172 56242 46228 56252
rect 41132 56130 41188 56140
rect 42140 56196 42196 56206
rect 42140 56102 42196 56140
rect 44940 56196 44996 56206
rect 41244 56082 41300 56094
rect 41244 56030 41246 56082
rect 41298 56030 41300 56082
rect 40348 55970 40404 55982
rect 40348 55918 40350 55970
rect 40402 55918 40404 55970
rect 40348 55412 40404 55918
rect 40348 54628 40404 55356
rect 41244 55412 41300 56030
rect 41244 55346 41300 55356
rect 42588 56084 42644 56094
rect 40348 54562 40404 54572
rect 39788 53902 39790 53954
rect 39842 53902 39844 53954
rect 39788 53890 39844 53902
rect 39228 53844 39284 53854
rect 39228 53750 39284 53788
rect 42364 53844 42420 53854
rect 42364 53750 42420 53788
rect 41580 53732 41636 53742
rect 38444 53678 38446 53730
rect 38498 53678 38500 53730
rect 38444 53666 38500 53678
rect 41244 53730 41636 53732
rect 41244 53678 41582 53730
rect 41634 53678 41636 53730
rect 41244 53676 41636 53678
rect 39116 53508 39172 53518
rect 39116 53414 39172 53452
rect 39564 53508 39620 53518
rect 39452 52836 39508 52846
rect 39564 52836 39620 53452
rect 39452 52834 39620 52836
rect 39452 52782 39454 52834
rect 39506 52782 39620 52834
rect 39452 52780 39620 52782
rect 39452 52770 39508 52780
rect 37548 51268 37604 51278
rect 36764 50484 36820 50494
rect 36092 50370 36148 50382
rect 36092 50318 36094 50370
rect 36146 50318 36148 50370
rect 36092 49812 36148 50318
rect 36652 50370 36708 50382
rect 36652 50318 36654 50370
rect 36706 50318 36708 50370
rect 36428 49812 36484 49822
rect 36652 49812 36708 50318
rect 36092 49810 36708 49812
rect 36092 49758 36430 49810
rect 36482 49758 36708 49810
rect 36092 49756 36708 49758
rect 35980 49644 36148 49700
rect 35868 49140 35924 49150
rect 35868 49046 35924 49084
rect 35756 48860 35924 48916
rect 33852 48692 33908 48702
rect 32956 46564 33012 46574
rect 32396 46002 32676 46004
rect 32396 45950 32398 46002
rect 32450 45950 32676 46002
rect 32396 45948 32676 45950
rect 32396 45938 32452 45948
rect 31724 45378 31780 45388
rect 32620 45330 32676 45948
rect 32620 45278 32622 45330
rect 32674 45278 32676 45330
rect 31612 44370 31668 44380
rect 31948 45220 32004 45230
rect 31948 44434 32004 45164
rect 32172 45220 32228 45230
rect 32172 45126 32228 45164
rect 32620 45220 32676 45278
rect 32620 45154 32676 45164
rect 32060 44882 32116 44894
rect 32060 44830 32062 44882
rect 32114 44830 32116 44882
rect 32060 44772 32116 44830
rect 32060 44706 32116 44716
rect 31948 44382 31950 44434
rect 32002 44382 32004 44434
rect 31948 44370 32004 44382
rect 32508 44210 32564 44222
rect 32508 44158 32510 44210
rect 32562 44158 32564 44210
rect 31836 44098 31892 44110
rect 31836 44046 31838 44098
rect 31890 44046 31892 44098
rect 31276 43586 31332 43596
rect 31612 43652 31668 43662
rect 31612 43558 31668 43596
rect 31500 43314 31556 43326
rect 31500 43262 31502 43314
rect 31554 43262 31556 43314
rect 31500 43092 31556 43262
rect 31500 43026 31556 43036
rect 31612 42196 31668 42206
rect 31388 42084 31444 42094
rect 31052 40628 31108 40638
rect 31052 40514 31108 40572
rect 31388 40626 31444 42028
rect 31388 40574 31390 40626
rect 31442 40574 31444 40626
rect 31388 40562 31444 40574
rect 31052 40462 31054 40514
rect 31106 40462 31108 40514
rect 31052 40450 31108 40462
rect 31164 40516 31220 40526
rect 31164 40422 31220 40460
rect 31276 39508 31332 39518
rect 30492 38210 30548 38220
rect 30604 38612 30772 38668
rect 30828 39340 30996 39396
rect 31052 39452 31276 39508
rect 30828 38668 30884 39340
rect 30940 39060 30996 39070
rect 31052 39060 31108 39452
rect 31276 39414 31332 39452
rect 31500 39506 31556 39518
rect 31500 39454 31502 39506
rect 31554 39454 31556 39506
rect 30996 39004 31108 39060
rect 30940 38928 30996 39004
rect 30828 38612 31332 38668
rect 30604 38052 30660 38612
rect 30492 37996 30660 38052
rect 30828 38052 30884 38062
rect 31164 38052 31220 38062
rect 30828 38050 31220 38052
rect 30828 37998 30830 38050
rect 30882 37998 31166 38050
rect 31218 37998 31220 38050
rect 30828 37996 31220 37998
rect 30156 37886 30158 37938
rect 30210 37886 30212 37938
rect 29932 35746 29988 35756
rect 29372 35252 29428 35262
rect 27916 34468 27972 34478
rect 27916 34020 27972 34412
rect 27132 33182 27134 33234
rect 27186 33182 27188 33234
rect 26796 33012 26852 33022
rect 26852 32956 26964 33012
rect 26796 32946 26852 32956
rect 26684 32510 26686 32562
rect 26738 32510 26740 32562
rect 26684 32498 26740 32510
rect 26908 32788 26964 32956
rect 26908 31890 26964 32732
rect 27132 32676 27188 33182
rect 27356 33180 27524 33236
rect 27804 33236 27860 33246
rect 27076 32620 27188 32676
rect 27244 32900 27300 32910
rect 27244 32786 27300 32844
rect 27244 32734 27246 32786
rect 27298 32734 27300 32786
rect 27244 32676 27300 32734
rect 27356 32786 27412 33180
rect 27692 33124 27748 33162
rect 27804 33142 27860 33180
rect 27692 33058 27748 33068
rect 27356 32734 27358 32786
rect 27410 32734 27412 32786
rect 27356 32722 27412 32734
rect 27468 33012 27524 33022
rect 27468 32786 27524 32956
rect 27916 32900 27972 33964
rect 28476 34468 28532 34478
rect 28476 33796 28532 34412
rect 28476 33730 28532 33740
rect 27468 32734 27470 32786
rect 27522 32734 27524 32786
rect 27468 32722 27524 32734
rect 27692 32844 27972 32900
rect 28028 33236 28084 33246
rect 27076 32228 27132 32620
rect 27244 32610 27300 32620
rect 27580 32676 27636 32686
rect 27580 32562 27636 32620
rect 27580 32510 27582 32562
rect 27634 32510 27636 32562
rect 27580 32498 27636 32510
rect 27692 32340 27748 32844
rect 27916 32340 27972 32350
rect 27356 32284 27748 32340
rect 27804 32338 27972 32340
rect 27804 32286 27918 32338
rect 27970 32286 27972 32338
rect 27804 32284 27972 32286
rect 27076 32172 27188 32228
rect 26908 31838 26910 31890
rect 26962 31838 26964 31890
rect 26908 31826 26964 31838
rect 26236 29538 26516 29540
rect 26236 29486 26238 29538
rect 26290 29486 26516 29538
rect 26236 29484 26516 29486
rect 26236 29474 26292 29484
rect 25340 27246 25342 27298
rect 25394 27246 25396 27298
rect 25340 27234 25396 27246
rect 25676 28980 25732 28990
rect 25228 26852 25284 26908
rect 24556 26450 24612 26460
rect 24108 25732 24164 25742
rect 23996 25730 24164 25732
rect 23996 25678 24110 25730
rect 24162 25678 24164 25730
rect 23996 25676 24164 25678
rect 24108 25666 24164 25676
rect 23996 25394 24052 25406
rect 23996 25342 23998 25394
rect 24050 25342 24052 25394
rect 23212 25004 23604 25060
rect 23212 24946 23268 25004
rect 23212 24894 23214 24946
rect 23266 24894 23268 24946
rect 23212 24882 23268 24894
rect 23548 24948 23604 25004
rect 22428 24770 22484 24780
rect 22428 24612 22484 24622
rect 22428 24518 22484 24556
rect 22764 24612 22820 24622
rect 22764 23938 22820 24556
rect 22764 23886 22766 23938
rect 22818 23886 22820 23938
rect 22092 23378 22260 23380
rect 22092 23326 22094 23378
rect 22146 23326 22260 23378
rect 22092 23324 22260 23326
rect 22316 23828 22372 23838
rect 22092 23314 22148 23324
rect 22316 23154 22372 23772
rect 22316 23102 22318 23154
rect 22370 23102 22372 23154
rect 22316 23090 22372 23102
rect 22764 23154 22820 23886
rect 23212 23828 23268 23838
rect 23212 23734 23268 23772
rect 23100 23716 23156 23726
rect 22988 23604 23044 23614
rect 22988 23266 23044 23548
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22988 23202 23044 23214
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 21980 22978 22036 22988
rect 22764 23044 22820 23102
rect 23100 23154 23156 23660
rect 23548 23604 23604 24892
rect 23660 25172 23716 25182
rect 23660 24612 23716 25116
rect 23996 24724 24052 25342
rect 24108 25284 24164 25294
rect 24108 25190 24164 25228
rect 24668 25282 24724 25294
rect 24668 25230 24670 25282
rect 24722 25230 24724 25282
rect 24668 25172 24724 25230
rect 24668 25106 24724 25116
rect 23996 24658 24052 24668
rect 24108 25060 24164 25070
rect 23660 24518 23716 24556
rect 23548 23378 23604 23548
rect 23548 23326 23550 23378
rect 23602 23326 23604 23378
rect 23548 23314 23604 23326
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 23100 23090 23156 23102
rect 22764 22978 22820 22988
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 12348 4498 12404 4508
rect 16492 5348 16548 5358
rect 16492 4562 16548 5292
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 16492 4510 16494 4562
rect 16546 4510 16548 4562
rect 15260 3668 15316 3678
rect 11788 3602 11844 3612
rect 14924 3666 15316 3668
rect 14924 3614 15262 3666
rect 15314 3614 15316 3666
rect 14924 3612 15316 3614
rect 10892 3554 11172 3556
rect 10892 3502 10894 3554
rect 10946 3502 11172 3554
rect 10892 3500 11172 3502
rect 10892 3490 10948 3500
rect 6076 3330 6356 3332
rect 6076 3278 6078 3330
rect 6130 3278 6356 3330
rect 6076 3276 6356 3278
rect 8876 3444 8932 3454
rect 6076 3266 6132 3276
rect 8876 800 8932 3388
rect 9996 3444 10052 3454
rect 9996 3350 10052 3388
rect 11676 3332 11732 3342
rect 11564 3330 11732 3332
rect 11564 3278 11678 3330
rect 11730 3278 11732 3330
rect 11564 3276 11732 3278
rect 11564 800 11620 3276
rect 11676 3266 11732 3276
rect 14924 800 14980 3612
rect 15260 3602 15316 3612
rect 16268 3556 16324 3566
rect 16492 3556 16548 4510
rect 16828 3668 16884 3678
rect 16828 3574 16884 3612
rect 17724 3668 17780 3678
rect 16268 3554 16548 3556
rect 16268 3502 16270 3554
rect 16322 3502 16548 3554
rect 16268 3500 16548 3502
rect 17724 3554 17780 3612
rect 17724 3502 17726 3554
rect 17778 3502 17780 3554
rect 16268 3490 16324 3500
rect 17724 3490 17780 3502
rect 18396 3666 18452 3678
rect 18396 3614 18398 3666
rect 18450 3614 18452 3666
rect 17612 812 17780 868
rect 17612 800 17668 812
rect 5292 728 5544 800
rect 5320 200 5544 728
rect 8680 728 8932 800
rect 11368 728 11620 800
rect 14728 728 14980 800
rect 17416 728 17668 800
rect 17724 756 17780 812
rect 18396 756 18452 3614
rect 20748 3444 20804 3454
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 8680 200 8904 728
rect 11368 200 11592 728
rect 14728 200 14952 728
rect 17416 200 17640 728
rect 17724 700 18452 756
rect 20748 800 20804 3388
rect 21420 3444 21476 3454
rect 21420 3350 21476 3388
rect 23324 3444 23380 3454
rect 23772 3444 23828 3454
rect 23324 3442 23828 3444
rect 23324 3390 23326 3442
rect 23378 3390 23774 3442
rect 23826 3390 23828 3442
rect 23324 3388 23828 3390
rect 23324 3378 23380 3388
rect 21756 3332 21812 3342
rect 21756 3238 21812 3276
rect 23548 800 23604 3388
rect 23772 3378 23828 3388
rect 24108 3330 24164 25004
rect 24332 24948 24388 24958
rect 24220 24724 24276 24734
rect 24220 24052 24276 24668
rect 24220 23986 24276 23996
rect 24332 24164 24388 24892
rect 24668 24948 24724 24958
rect 24668 24854 24724 24892
rect 24780 24948 24836 24958
rect 24892 24948 24948 26852
rect 24780 24946 24948 24948
rect 24780 24894 24782 24946
rect 24834 24894 24948 24946
rect 24780 24892 24948 24894
rect 25116 26796 25284 26852
rect 25676 27188 25732 28924
rect 26460 28980 26516 29484
rect 26460 28914 26516 28924
rect 26908 30100 26964 30110
rect 26460 28756 26516 28766
rect 26460 28662 26516 28700
rect 26908 28756 26964 30044
rect 26908 28690 26964 28700
rect 27020 28532 27076 28542
rect 26908 28530 27076 28532
rect 26908 28478 27022 28530
rect 27074 28478 27076 28530
rect 26908 28476 27076 28478
rect 24780 24882 24836 24892
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24444 24612 24500 24670
rect 24444 24546 24500 24556
rect 24332 23938 24388 24108
rect 25116 24050 25172 26796
rect 25676 26514 25732 27132
rect 26012 27300 26068 27310
rect 26012 27186 26068 27244
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27122 26068 27134
rect 26460 26964 26516 27002
rect 26460 26898 26516 26908
rect 25676 26462 25678 26514
rect 25730 26462 25732 26514
rect 25676 26450 25732 26462
rect 26908 26404 26964 28476
rect 27020 28466 27076 28476
rect 27132 27524 27188 32172
rect 27244 32116 27300 32126
rect 27244 31890 27300 32060
rect 27244 31838 27246 31890
rect 27298 31838 27300 31890
rect 27244 31826 27300 31838
rect 27132 27458 27188 27468
rect 27020 27300 27076 27310
rect 27020 26962 27076 27244
rect 27020 26910 27022 26962
rect 27074 26910 27076 26962
rect 27020 26898 27076 26910
rect 27356 26908 27412 32284
rect 27468 28756 27524 28766
rect 27468 28642 27524 28700
rect 27468 28590 27470 28642
rect 27522 28590 27524 28642
rect 27468 28578 27524 28590
rect 27692 27076 27748 27114
rect 27692 27010 27748 27020
rect 27804 26908 27860 32284
rect 27916 32274 27972 32284
rect 28028 30100 28084 33180
rect 28252 33236 28308 33246
rect 28252 33142 28308 33180
rect 28924 33236 28980 33246
rect 28924 33122 28980 33180
rect 28924 33070 28926 33122
rect 28978 33070 28980 33122
rect 28588 32900 28644 32910
rect 28588 32786 28644 32844
rect 28588 32734 28590 32786
rect 28642 32734 28644 32786
rect 28588 32722 28644 32734
rect 28924 32564 28980 33070
rect 28924 32498 28980 32508
rect 28140 32338 28196 32350
rect 28140 32286 28142 32338
rect 28194 32286 28196 32338
rect 28140 31892 28196 32286
rect 29372 32340 29428 35196
rect 30156 35252 30212 37886
rect 30380 37940 30436 37950
rect 30380 37846 30436 37884
rect 30492 36594 30548 37996
rect 30828 37986 30884 37996
rect 31164 37986 31220 37996
rect 30604 37828 30660 37838
rect 30604 37826 31108 37828
rect 30604 37774 30606 37826
rect 30658 37774 31108 37826
rect 30604 37772 31108 37774
rect 30604 37762 30660 37772
rect 30940 37380 30996 37390
rect 30940 37286 30996 37324
rect 31052 36706 31108 37772
rect 31276 37380 31332 38612
rect 31500 38052 31556 39454
rect 31612 39394 31668 42140
rect 31724 40964 31780 40974
rect 31724 39620 31780 40908
rect 31836 40516 31892 44046
rect 32508 43762 32564 44158
rect 32508 43710 32510 43762
rect 32562 43710 32564 43762
rect 32060 43652 32116 43662
rect 32060 43558 32116 43596
rect 32396 43316 32452 43326
rect 32060 40628 32116 40638
rect 31836 40450 31892 40460
rect 31948 40572 32060 40628
rect 31836 40292 31892 40302
rect 31836 40198 31892 40236
rect 31836 39620 31892 39630
rect 31724 39618 31892 39620
rect 31724 39566 31838 39618
rect 31890 39566 31892 39618
rect 31724 39564 31892 39566
rect 31836 39554 31892 39564
rect 31612 39342 31614 39394
rect 31666 39342 31668 39394
rect 31612 39330 31668 39342
rect 31948 38948 32004 40572
rect 32060 40534 32116 40572
rect 31948 38882 32004 38892
rect 32060 40290 32116 40302
rect 32060 40238 32062 40290
rect 32114 40238 32116 40290
rect 31500 37958 31556 37996
rect 31948 37940 32004 37950
rect 31276 37314 31332 37324
rect 31388 37826 31444 37838
rect 31388 37774 31390 37826
rect 31442 37774 31444 37826
rect 31052 36654 31054 36706
rect 31106 36654 31108 36706
rect 31052 36642 31108 36654
rect 30492 36542 30494 36594
rect 30546 36542 30548 36594
rect 30492 36530 30548 36542
rect 30604 36484 30660 36494
rect 30604 36390 30660 36428
rect 30716 36482 30772 36494
rect 30716 36430 30718 36482
rect 30770 36430 30772 36482
rect 30380 36260 30436 36270
rect 30380 36166 30436 36204
rect 30716 35812 30772 36430
rect 30716 35746 30772 35756
rect 31276 36482 31332 36494
rect 31276 36430 31278 36482
rect 31330 36430 31332 36482
rect 31276 35588 31332 36430
rect 31388 36484 31444 37774
rect 31948 37826 32004 37884
rect 31948 37774 31950 37826
rect 32002 37774 32004 37826
rect 31500 37380 31556 37390
rect 31500 37286 31556 37324
rect 31948 37156 32004 37774
rect 32060 37492 32116 40238
rect 32284 39508 32340 39518
rect 32284 39414 32340 39452
rect 32060 37426 32116 37436
rect 32396 37828 32452 43260
rect 32508 38164 32564 43710
rect 32620 44098 32676 44110
rect 32620 44046 32622 44098
rect 32674 44046 32676 44098
rect 32620 43428 32676 44046
rect 32620 43362 32676 43372
rect 32956 43316 33012 46508
rect 33740 46564 33796 46574
rect 33740 46470 33796 46508
rect 33628 46450 33684 46462
rect 33628 46398 33630 46450
rect 33682 46398 33684 46450
rect 33628 45332 33684 46398
rect 33516 44436 33572 44446
rect 33068 44098 33124 44110
rect 33068 44046 33070 44098
rect 33122 44046 33124 44098
rect 33068 43652 33124 44046
rect 33516 43708 33572 44380
rect 33628 44324 33684 45276
rect 33628 44258 33684 44268
rect 33516 43652 33684 43708
rect 33068 43586 33124 43596
rect 33628 43428 33684 43652
rect 33852 43652 33908 48636
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34412 46564 34468 46574
rect 34860 46564 34916 46574
rect 34412 46562 34916 46564
rect 34412 46510 34414 46562
rect 34466 46510 34862 46562
rect 34914 46510 34916 46562
rect 34412 46508 34916 46510
rect 34412 46498 34468 46508
rect 34300 46450 34356 46462
rect 34300 46398 34302 46450
rect 34354 46398 34356 46450
rect 34076 45780 34132 45790
rect 34076 45686 34132 45724
rect 33964 45666 34020 45678
rect 33964 45614 33966 45666
rect 34018 45614 34020 45666
rect 33964 44212 34020 45614
rect 33964 44146 34020 44156
rect 34076 44324 34132 44334
rect 33964 43652 34020 43662
rect 33852 43650 34020 43652
rect 33852 43598 33966 43650
rect 34018 43598 34020 43650
rect 33852 43596 34020 43598
rect 33964 43586 34020 43596
rect 33852 43428 33908 43438
rect 33628 43426 33908 43428
rect 33628 43374 33854 43426
rect 33906 43374 33908 43426
rect 33628 43372 33908 43374
rect 33852 43362 33908 43372
rect 32956 43250 33012 43260
rect 33740 42754 33796 42766
rect 33740 42702 33742 42754
rect 33794 42702 33796 42754
rect 33740 42084 33796 42702
rect 33740 42018 33796 42028
rect 32620 41748 32676 41758
rect 32620 40628 32676 41692
rect 34076 41300 34132 44268
rect 34188 43652 34244 43662
rect 34188 43428 34244 43596
rect 34300 43540 34356 46398
rect 34524 45780 34580 46508
rect 34860 46498 34916 46508
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35868 46114 35924 48860
rect 35868 46062 35870 46114
rect 35922 46062 35924 46114
rect 35420 46002 35476 46014
rect 35420 45950 35422 46002
rect 35474 45950 35476 46002
rect 35420 45892 35476 45950
rect 35532 45892 35588 45902
rect 35420 45890 35588 45892
rect 35420 45838 35534 45890
rect 35586 45838 35588 45890
rect 35420 45836 35588 45838
rect 35532 45826 35588 45836
rect 35644 45892 35700 45902
rect 34524 45686 34580 45724
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34300 43474 34356 43484
rect 35084 43540 35140 43550
rect 35084 43538 35252 43540
rect 35084 43486 35086 43538
rect 35138 43486 35252 43538
rect 35084 43484 35252 43486
rect 35084 43474 35140 43484
rect 35196 43428 35252 43484
rect 35532 43428 35588 43438
rect 35196 43426 35588 43428
rect 35196 43374 35534 43426
rect 35586 43374 35588 43426
rect 35196 43372 35588 43374
rect 34188 42754 34244 43372
rect 34748 43314 34804 43326
rect 34748 43262 34750 43314
rect 34802 43262 34804 43314
rect 34636 42868 34692 42878
rect 34748 42868 34804 43262
rect 35084 43316 35140 43326
rect 35084 43222 35140 43260
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34636 42866 34804 42868
rect 34636 42814 34638 42866
rect 34690 42814 34804 42866
rect 34636 42812 34804 42814
rect 34636 42802 34692 42812
rect 34188 42702 34190 42754
rect 34242 42702 34244 42754
rect 34188 42690 34244 42702
rect 35532 42084 35588 43372
rect 35420 42028 35588 42084
rect 35420 41748 35476 42028
rect 35420 41682 35476 41692
rect 35532 41860 35588 41870
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41412 35588 41804
rect 35644 41524 35700 45836
rect 35756 45892 35812 45902
rect 35868 45892 35924 46062
rect 35756 45890 35924 45892
rect 35756 45838 35758 45890
rect 35810 45838 35924 45890
rect 35756 45836 35924 45838
rect 35756 45826 35812 45836
rect 35980 45666 36036 45678
rect 35980 45614 35982 45666
rect 36034 45614 36036 45666
rect 35980 45556 36036 45614
rect 35980 45490 36036 45500
rect 36092 43708 36148 49644
rect 36428 48804 36484 49756
rect 36764 49700 36820 50428
rect 36428 48710 36484 48748
rect 36652 49644 36820 49700
rect 36876 49700 36932 49710
rect 36876 49698 37044 49700
rect 36876 49646 36878 49698
rect 36930 49646 37044 49698
rect 36876 49644 37044 49646
rect 36204 45890 36260 45902
rect 36204 45838 36206 45890
rect 36258 45838 36260 45890
rect 36204 45668 36260 45838
rect 36652 45892 36708 49644
rect 36876 49634 36932 49644
rect 36988 48804 37044 49644
rect 36652 45826 36708 45836
rect 36764 48356 36820 48366
rect 36652 45668 36708 45678
rect 36204 45666 36708 45668
rect 36204 45614 36654 45666
rect 36706 45614 36708 45666
rect 36204 45612 36708 45614
rect 36652 44996 36708 45612
rect 36652 44930 36708 44940
rect 35644 41458 35700 41468
rect 35868 43652 36148 43708
rect 36764 43762 36820 48300
rect 36988 45780 37044 48748
rect 37436 48804 37492 48814
rect 37436 48710 37492 48748
rect 37100 46562 37156 46574
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 37100 45892 37156 46510
rect 37100 45826 37156 45836
rect 37436 46564 37492 46574
rect 37548 46564 37604 51212
rect 38556 51268 38612 51278
rect 38556 51174 38612 51212
rect 39004 51266 39060 51278
rect 39004 51214 39006 51266
rect 39058 51214 39060 51266
rect 39004 50820 39060 51214
rect 39452 51044 39508 51054
rect 39116 50820 39172 50830
rect 39004 50818 39172 50820
rect 39004 50766 39118 50818
rect 39170 50766 39172 50818
rect 39004 50764 39172 50766
rect 37436 46562 37604 46564
rect 37436 46510 37438 46562
rect 37490 46510 37604 46562
rect 37436 46508 37604 46510
rect 37772 49812 37828 49822
rect 36988 45714 37044 45724
rect 37436 45668 37492 46508
rect 37660 45668 37716 45678
rect 37436 45666 37716 45668
rect 37436 45614 37662 45666
rect 37714 45614 37716 45666
rect 37436 45612 37716 45614
rect 37324 45220 37380 45230
rect 37324 45126 37380 45164
rect 36764 43710 36766 43762
rect 36818 43710 36820 43762
rect 36764 43698 36820 43710
rect 36988 45106 37044 45118
rect 36988 45054 36990 45106
rect 37042 45054 37044 45106
rect 36988 44996 37044 45054
rect 36876 43652 36932 43662
rect 34188 41300 34244 41310
rect 33628 41298 34244 41300
rect 33628 41246 34190 41298
rect 34242 41246 34244 41298
rect 33628 41244 34244 41246
rect 33628 41074 33684 41244
rect 34188 41234 34244 41244
rect 35308 41300 35364 41310
rect 33628 41022 33630 41074
rect 33682 41022 33684 41074
rect 33628 41010 33684 41022
rect 33740 41074 33796 41086
rect 33740 41022 33742 41074
rect 33794 41022 33796 41074
rect 33404 40964 33460 40974
rect 33404 40870 33460 40908
rect 32620 40496 32676 40572
rect 32508 38098 32564 38108
rect 33068 40292 33124 40302
rect 32844 38052 32900 38062
rect 32844 37958 32900 37996
rect 32956 37828 33012 37838
rect 32396 37826 33012 37828
rect 32396 37774 32398 37826
rect 32450 37774 32958 37826
rect 33010 37774 33012 37826
rect 32396 37772 33012 37774
rect 31948 37090 32004 37100
rect 32284 36820 32340 36830
rect 32284 36594 32340 36764
rect 32284 36542 32286 36594
rect 32338 36542 32340 36594
rect 32284 36530 32340 36542
rect 31388 36418 31444 36428
rect 32172 36484 32228 36494
rect 32172 36390 32228 36428
rect 32396 35700 32452 37772
rect 32956 37762 33012 37772
rect 32620 37492 32676 37502
rect 32620 37398 32676 37436
rect 32732 36820 32788 36830
rect 32732 36594 32788 36764
rect 32732 36542 32734 36594
rect 32786 36542 32788 36594
rect 32732 35924 32788 36542
rect 32844 35924 32900 35934
rect 32732 35922 32900 35924
rect 32732 35870 32846 35922
rect 32898 35870 32900 35922
rect 32732 35868 32900 35870
rect 32396 35606 32452 35644
rect 31500 35588 31556 35598
rect 31276 35586 31556 35588
rect 31276 35534 31502 35586
rect 31554 35534 31556 35586
rect 31276 35532 31556 35534
rect 31500 35476 31556 35532
rect 32844 35588 32900 35868
rect 32844 35522 32900 35532
rect 31500 35410 31556 35420
rect 30156 35186 30212 35196
rect 29596 35140 29652 35150
rect 29596 35046 29652 35084
rect 29708 34802 29764 34814
rect 29708 34750 29710 34802
rect 29762 34750 29764 34802
rect 29708 34692 29764 34750
rect 30156 34692 30212 34702
rect 29708 34690 30212 34692
rect 29708 34638 30158 34690
rect 30210 34638 30212 34690
rect 29708 34636 30212 34638
rect 29484 34580 29540 34590
rect 29484 33460 29540 34524
rect 29708 34132 29764 34636
rect 30156 34626 30212 34636
rect 29708 34066 29764 34076
rect 32620 33572 32676 33582
rect 33068 33572 33124 40236
rect 33180 40068 33236 40078
rect 33180 39394 33236 40012
rect 33740 39732 33796 41022
rect 35084 41076 35140 41086
rect 34636 40964 34692 40974
rect 33852 40404 33908 40414
rect 33852 39842 33908 40348
rect 34300 40402 34356 40414
rect 34300 40350 34302 40402
rect 34354 40350 34356 40402
rect 34300 40292 34356 40350
rect 34300 40226 34356 40236
rect 33852 39790 33854 39842
rect 33906 39790 33908 39842
rect 33852 39778 33908 39790
rect 34076 40180 34132 40190
rect 33180 39342 33182 39394
rect 33234 39342 33236 39394
rect 33180 39284 33236 39342
rect 33180 39218 33236 39228
rect 33628 39676 33796 39732
rect 33516 38050 33572 38062
rect 33516 37998 33518 38050
rect 33570 37998 33572 38050
rect 33180 37826 33236 37838
rect 33180 37774 33182 37826
rect 33234 37774 33236 37826
rect 33180 37492 33236 37774
rect 33180 37044 33236 37436
rect 33180 35812 33236 36988
rect 33516 36708 33572 37998
rect 33516 36642 33572 36652
rect 33516 36484 33572 36494
rect 33516 36390 33572 36428
rect 33628 36036 33684 39676
rect 33740 39506 33796 39518
rect 33740 39454 33742 39506
rect 33794 39454 33796 39506
rect 33740 39284 33796 39454
rect 33740 39218 33796 39228
rect 33964 38052 34020 38062
rect 33964 37268 34020 37996
rect 33964 37202 34020 37212
rect 34076 36932 34132 40124
rect 34524 39956 34580 39966
rect 34524 39396 34580 39900
rect 34636 39844 34692 40908
rect 35084 40962 35140 41020
rect 35084 40910 35086 40962
rect 35138 40910 35140 40962
rect 34860 40628 34916 40638
rect 34860 40534 34916 40572
rect 35084 40516 35140 40910
rect 35084 40450 35140 40460
rect 34972 40404 35028 40414
rect 34748 40180 34804 40190
rect 34748 40086 34804 40124
rect 34636 39778 34692 39788
rect 34524 39330 34580 39340
rect 34748 39506 34804 39518
rect 34748 39454 34750 39506
rect 34802 39454 34804 39506
rect 34412 38724 34468 38734
rect 34748 38724 34804 39454
rect 34860 39508 34916 39518
rect 34972 39508 35028 40348
rect 35084 40292 35140 40302
rect 35308 40292 35364 41244
rect 35532 41300 35588 41356
rect 35532 41298 35812 41300
rect 35532 41246 35534 41298
rect 35586 41246 35812 41298
rect 35532 41244 35812 41246
rect 35532 41234 35588 41244
rect 35756 40626 35812 41244
rect 35756 40574 35758 40626
rect 35810 40574 35812 40626
rect 35756 40562 35812 40574
rect 35868 40626 35924 43652
rect 36876 43558 36932 43596
rect 36652 43540 36708 43550
rect 35980 43428 36036 43438
rect 35980 43334 36036 43372
rect 36204 42532 36260 42542
rect 36204 42438 36260 42476
rect 36652 42532 36708 43484
rect 36988 43316 37044 44940
rect 37212 44994 37268 45006
rect 37212 44942 37214 44994
rect 37266 44942 37268 44994
rect 36652 42466 36708 42476
rect 36764 43260 37044 43316
rect 37100 43428 37156 43438
rect 36428 41300 36484 41310
rect 36428 41206 36484 41244
rect 35868 40574 35870 40626
rect 35922 40574 35924 40626
rect 35868 40562 35924 40574
rect 35980 41076 36036 41086
rect 35980 40628 36036 41020
rect 35980 40562 36036 40572
rect 36204 40516 36260 40526
rect 35980 40404 36036 40414
rect 35980 40310 36036 40348
rect 36204 40402 36260 40460
rect 36204 40350 36206 40402
rect 36258 40350 36260 40402
rect 36204 40338 36260 40350
rect 36540 40404 36596 40414
rect 35084 40290 35364 40292
rect 35084 40238 35086 40290
rect 35138 40238 35364 40290
rect 35084 40236 35364 40238
rect 35084 40226 35140 40236
rect 36428 40178 36484 40190
rect 36428 40126 36430 40178
rect 36482 40126 36484 40178
rect 35644 40068 35700 40078
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39620 35140 39630
rect 35084 39526 35140 39564
rect 35644 39618 35700 40012
rect 36428 39732 36484 40126
rect 36428 39666 36484 39676
rect 35644 39566 35646 39618
rect 35698 39566 35700 39618
rect 34860 39506 35028 39508
rect 34860 39454 34862 39506
rect 34914 39454 35028 39506
rect 34860 39452 35028 39454
rect 34860 39442 34916 39452
rect 35084 39396 35140 39406
rect 34972 39060 35028 39070
rect 35084 39060 35140 39340
rect 35644 39284 35700 39566
rect 36204 39506 36260 39518
rect 36204 39454 36206 39506
rect 36258 39454 36260 39506
rect 35756 39396 35812 39434
rect 35980 39396 36036 39406
rect 35756 39330 35812 39340
rect 35868 39394 36036 39396
rect 35868 39342 35982 39394
rect 36034 39342 36036 39394
rect 35868 39340 36036 39342
rect 34972 39058 35140 39060
rect 34972 39006 34974 39058
rect 35026 39006 35140 39058
rect 34972 39004 35140 39006
rect 35420 39060 35476 39070
rect 35644 39060 35700 39228
rect 35420 39058 35700 39060
rect 35420 39006 35422 39058
rect 35474 39006 35700 39058
rect 35420 39004 35700 39006
rect 35756 39172 35812 39182
rect 35756 39058 35812 39116
rect 35756 39006 35758 39058
rect 35810 39006 35812 39058
rect 34972 38994 35028 39004
rect 35420 38994 35476 39004
rect 35756 38994 35812 39006
rect 33628 35970 33684 35980
rect 33964 36876 34132 36932
rect 34188 38722 34804 38724
rect 34188 38670 34414 38722
rect 34466 38670 34804 38722
rect 34188 38668 34804 38670
rect 33628 35812 33684 35822
rect 33236 35756 33348 35812
rect 33180 35746 33236 35756
rect 33292 35026 33348 35756
rect 33964 35812 34020 36876
rect 34076 36708 34132 36718
rect 34076 36614 34132 36652
rect 34076 36484 34132 36494
rect 34188 36484 34244 38668
rect 34412 38658 34468 38668
rect 35868 38612 35924 39340
rect 35980 39330 36036 39340
rect 36204 39172 36260 39454
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34412 38164 34468 38174
rect 34412 38070 34468 38108
rect 35084 38164 35140 38174
rect 35084 38070 35140 38108
rect 35308 38052 35364 38062
rect 35308 37958 35364 37996
rect 35084 37156 35140 37166
rect 34972 36708 35028 36718
rect 34412 36596 34468 36606
rect 34132 36428 34244 36484
rect 34300 36540 34412 36596
rect 34076 36390 34132 36428
rect 33964 35756 34132 35812
rect 33628 35718 33684 35756
rect 33740 35698 33796 35710
rect 33740 35646 33742 35698
rect 33794 35646 33796 35698
rect 33740 35588 33796 35646
rect 33740 35308 33796 35532
rect 33740 35252 34020 35308
rect 33292 34974 33294 35026
rect 33346 34974 33348 35026
rect 33292 34962 33348 34974
rect 33852 34132 33908 34142
rect 33852 34020 33908 34076
rect 32620 33570 33124 33572
rect 32620 33518 32622 33570
rect 32674 33518 33124 33570
rect 32620 33516 33124 33518
rect 33628 34018 33908 34020
rect 33628 33966 33854 34018
rect 33906 33966 33908 34018
rect 33628 33964 33908 33966
rect 32620 33506 32676 33516
rect 29708 33460 29764 33470
rect 29484 33404 29708 33460
rect 29596 33236 29652 33246
rect 29596 33142 29652 33180
rect 29708 33234 29764 33404
rect 30268 33460 30324 33470
rect 30268 33366 30324 33404
rect 29708 33182 29710 33234
rect 29762 33182 29764 33234
rect 29708 33170 29764 33182
rect 32284 33234 32340 33246
rect 32284 33182 32286 33234
rect 32338 33182 32340 33234
rect 29932 33122 29988 33134
rect 29932 33070 29934 33122
rect 29986 33070 29988 33122
rect 29372 32274 29428 32284
rect 29484 33012 29540 33022
rect 28140 31826 28196 31836
rect 29484 31220 29540 32956
rect 29932 31780 29988 33070
rect 31724 33124 31780 33134
rect 32284 33124 32340 33182
rect 31724 33122 32340 33124
rect 31724 33070 31726 33122
rect 31778 33070 32340 33122
rect 31724 33068 32340 33070
rect 32508 33122 32564 33134
rect 32508 33070 32510 33122
rect 32562 33070 32564 33122
rect 31724 33058 31780 33068
rect 30492 31892 30548 31902
rect 30492 31798 30548 31836
rect 29932 31714 29988 31724
rect 30828 31666 30884 31678
rect 30828 31614 30830 31666
rect 30882 31614 30884 31666
rect 30604 31554 30660 31566
rect 30604 31502 30606 31554
rect 30658 31502 30660 31554
rect 30604 31444 30660 31502
rect 30604 31378 30660 31388
rect 28924 31218 29540 31220
rect 28924 31166 29486 31218
rect 29538 31166 29540 31218
rect 28924 31164 29540 31166
rect 28924 30994 28980 31164
rect 29484 31154 29540 31164
rect 30828 31220 30884 31614
rect 30828 31154 30884 31164
rect 31276 31554 31332 31566
rect 31276 31502 31278 31554
rect 31330 31502 31332 31554
rect 31276 31220 31332 31502
rect 31724 31554 31780 31566
rect 31724 31502 31726 31554
rect 31778 31502 31780 31554
rect 31724 31444 31780 31502
rect 31724 31378 31780 31388
rect 31276 31154 31332 31164
rect 28924 30942 28926 30994
rect 28978 30942 28980 30994
rect 28924 30930 28980 30942
rect 28028 30034 28084 30044
rect 28140 30882 28196 30894
rect 28140 30830 28142 30882
rect 28194 30830 28196 30882
rect 28140 30772 28196 30830
rect 28700 30884 28756 30894
rect 28700 30790 28756 30828
rect 28588 30772 28644 30782
rect 28140 30770 28644 30772
rect 28140 30718 28590 30770
rect 28642 30718 28644 30770
rect 28140 30716 28644 30718
rect 28028 28868 28084 28878
rect 27916 28756 27972 28766
rect 27916 28662 27972 28700
rect 28028 28644 28084 28812
rect 27132 26852 27188 26862
rect 27020 26404 27076 26414
rect 26908 26402 27076 26404
rect 26908 26350 27022 26402
rect 27074 26350 27076 26402
rect 26908 26348 27076 26350
rect 27020 26338 27076 26348
rect 26908 25060 26964 25070
rect 26908 24946 26964 25004
rect 27132 25060 27188 26796
rect 27244 26852 27412 26908
rect 27468 26852 27860 26908
rect 27916 27748 27972 27758
rect 27916 27188 27972 27692
rect 27244 26516 27300 26852
rect 27244 26384 27300 26460
rect 27356 26180 27412 26190
rect 27468 26180 27524 26852
rect 27804 26516 27860 26526
rect 27804 26422 27860 26460
rect 27356 26178 27524 26180
rect 27356 26126 27358 26178
rect 27410 26126 27524 26178
rect 27356 26124 27524 26126
rect 27356 26114 27412 26124
rect 27132 24994 27188 25004
rect 26908 24894 26910 24946
rect 26962 24894 26964 24946
rect 26908 24882 26964 24894
rect 27468 24948 27524 24958
rect 27468 24854 27524 24892
rect 27804 24948 27860 24958
rect 27916 24948 27972 27132
rect 28028 27074 28084 28588
rect 28028 27022 28030 27074
rect 28082 27022 28084 27074
rect 28028 27010 28084 27022
rect 27804 24946 27972 24948
rect 27804 24894 27806 24946
rect 27858 24894 27972 24946
rect 27804 24892 27972 24894
rect 27804 24882 27860 24892
rect 27916 24836 27972 24892
rect 27916 24770 27972 24780
rect 25116 23998 25118 24050
rect 25170 23998 25172 24050
rect 25116 23986 25172 23998
rect 26348 24164 26404 24174
rect 26348 24050 26404 24108
rect 26348 23998 26350 24050
rect 26402 23998 26404 24050
rect 26348 23986 26404 23998
rect 24332 23886 24334 23938
rect 24386 23886 24388 23938
rect 24332 23874 24388 23886
rect 24220 23826 24276 23838
rect 24220 23774 24222 23826
rect 24274 23774 24276 23826
rect 24220 23716 24276 23774
rect 24220 23650 24276 23660
rect 27132 3332 27188 3342
rect 24108 3278 24110 3330
rect 24162 3278 24164 3330
rect 24108 3266 24164 3278
rect 27020 3330 27188 3332
rect 27020 3278 27134 3330
rect 27186 3278 27188 3330
rect 27020 3276 27188 3278
rect 27020 800 27076 3276
rect 27132 3266 27188 3276
rect 28140 3332 28196 30716
rect 28588 30706 28644 30716
rect 31164 29986 31220 29998
rect 31164 29934 31166 29986
rect 31218 29934 31220 29986
rect 28924 29316 28980 29326
rect 28476 29204 28532 29214
rect 28476 28756 28532 29148
rect 28252 27076 28308 27086
rect 28252 24946 28308 27020
rect 28476 26850 28532 28700
rect 28812 28756 28868 28766
rect 28588 28532 28644 28542
rect 28588 27300 28644 28476
rect 28700 28084 28756 28094
rect 28700 27990 28756 28028
rect 28812 27970 28868 28700
rect 28812 27918 28814 27970
rect 28866 27918 28868 27970
rect 28812 27906 28868 27918
rect 28700 27636 28756 27646
rect 28700 27542 28756 27580
rect 28588 26962 28644 27244
rect 28588 26910 28590 26962
rect 28642 26910 28644 26962
rect 28588 26898 28644 26910
rect 28700 27076 28756 27086
rect 28476 26798 28478 26850
rect 28530 26798 28532 26850
rect 28476 26786 28532 26798
rect 28252 24894 28254 24946
rect 28306 24894 28308 24946
rect 28252 24882 28308 24894
rect 28364 25060 28420 25070
rect 28364 24946 28420 25004
rect 28364 24894 28366 24946
rect 28418 24894 28420 24946
rect 28364 24882 28420 24894
rect 28588 24948 28644 24958
rect 28700 24948 28756 27020
rect 28924 25060 28980 29260
rect 29260 28532 29316 28542
rect 29260 28084 29316 28476
rect 31164 28532 31220 29934
rect 31164 28466 31220 28476
rect 31612 29988 31668 29998
rect 29260 27952 29316 28028
rect 29484 27300 29540 27310
rect 29484 27186 29540 27244
rect 29484 27134 29486 27186
rect 29538 27134 29540 27186
rect 29484 27122 29540 27134
rect 31276 27188 31332 27198
rect 31276 27094 31332 27132
rect 31612 27188 31668 29932
rect 31612 27122 31668 27132
rect 31724 27076 31780 27086
rect 31724 26982 31780 27020
rect 28924 24994 28980 25004
rect 28644 24892 28756 24948
rect 28588 24816 28644 24892
rect 28812 24836 28868 24846
rect 28812 11172 28868 24780
rect 28812 11106 28868 11116
rect 31836 8428 31892 33068
rect 32508 33012 32564 33070
rect 32508 32946 32564 32956
rect 33068 33122 33124 33134
rect 33068 33070 33070 33122
rect 33122 33070 33124 33122
rect 33068 33012 33124 33070
rect 33068 32946 33124 32956
rect 32060 32452 32116 32462
rect 32060 30434 32116 32396
rect 32060 30382 32062 30434
rect 32114 30382 32116 30434
rect 32060 30370 32116 30382
rect 33628 30212 33684 33964
rect 33852 33954 33908 33964
rect 33964 32788 34020 35252
rect 34076 33572 34132 35756
rect 34076 33506 34132 33516
rect 34188 35700 34244 35710
rect 33964 32656 34020 32732
rect 34188 32564 34244 35644
rect 34300 34356 34356 36540
rect 34412 36502 34468 36540
rect 34860 36596 34916 36606
rect 34860 36502 34916 36540
rect 34636 36484 34692 36494
rect 34412 35700 34468 35710
rect 34412 35606 34468 35644
rect 34524 34914 34580 34926
rect 34524 34862 34526 34914
rect 34578 34862 34580 34914
rect 34412 34356 34468 34366
rect 34300 34354 34468 34356
rect 34300 34302 34414 34354
rect 34466 34302 34468 34354
rect 34300 34300 34468 34302
rect 34412 33796 34468 34300
rect 34524 34354 34580 34862
rect 34524 34302 34526 34354
rect 34578 34302 34580 34354
rect 34524 34290 34580 34302
rect 34636 34132 34692 36428
rect 34860 36036 34916 36046
rect 34860 34914 34916 35980
rect 34972 35812 35028 36652
rect 34972 35698 35028 35756
rect 35084 35810 35140 37100
rect 35868 37044 35924 38556
rect 36092 38724 36148 38734
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 35758 35086 35810
rect 35138 35758 35140 35810
rect 35084 35746 35140 35758
rect 35532 36596 35588 36606
rect 34972 35646 34974 35698
rect 35026 35646 35028 35698
rect 34972 35634 35028 35646
rect 35196 35308 35460 35318
rect 34860 34862 34862 34914
rect 34914 34862 34916 34914
rect 34860 34850 34916 34862
rect 34972 35252 35028 35262
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34972 34916 35028 35196
rect 35532 35028 35588 36540
rect 35644 35812 35700 35822
rect 35644 35718 35700 35756
rect 35756 35812 35812 35822
rect 35868 35812 35924 36988
rect 35980 37938 36036 37950
rect 35980 37886 35982 37938
rect 36034 37886 36036 37938
rect 35980 36484 36036 37886
rect 35980 36418 36036 36428
rect 35980 36036 36036 36046
rect 35980 35922 36036 35980
rect 35980 35870 35982 35922
rect 36034 35870 36036 35922
rect 35980 35858 36036 35870
rect 35756 35810 35924 35812
rect 35756 35758 35758 35810
rect 35810 35758 35924 35810
rect 35756 35756 35924 35758
rect 35756 35746 35812 35756
rect 35756 35588 35812 35598
rect 35644 35028 35700 35038
rect 35532 35026 35700 35028
rect 35532 34974 35646 35026
rect 35698 34974 35700 35026
rect 35532 34972 35700 34974
rect 35644 34962 35700 34972
rect 35084 34916 35140 34926
rect 34972 34914 35140 34916
rect 34972 34862 35086 34914
rect 35138 34862 35140 34914
rect 34972 34860 35140 34862
rect 34636 34038 34692 34076
rect 34860 34690 34916 34702
rect 34860 34638 34862 34690
rect 34914 34638 34916 34690
rect 34412 33740 34804 33796
rect 34748 33570 34804 33740
rect 34748 33518 34750 33570
rect 34802 33518 34804 33570
rect 34748 33506 34804 33518
rect 34860 33572 34916 34638
rect 35084 34692 35140 34860
rect 35084 34626 35140 34636
rect 34860 33506 34916 33516
rect 34972 34356 35028 34366
rect 34972 33570 35028 34300
rect 34972 33518 34974 33570
rect 35026 33518 35028 33570
rect 34300 33124 34356 33134
rect 34300 33122 34692 33124
rect 34300 33070 34302 33122
rect 34354 33070 34692 33122
rect 34300 33068 34692 33070
rect 34300 33058 34356 33068
rect 34524 32788 34580 32798
rect 34524 32694 34580 32732
rect 34412 32564 34468 32574
rect 34188 32562 34468 32564
rect 34188 32510 34414 32562
rect 34466 32510 34468 32562
rect 34188 32508 34468 32510
rect 34076 31554 34132 31566
rect 34076 31502 34078 31554
rect 34130 31502 34132 31554
rect 34076 31444 34132 31502
rect 34300 31444 34356 32508
rect 34412 32498 34468 32508
rect 34076 31388 34356 31444
rect 32620 30098 32676 30110
rect 32620 30046 32622 30098
rect 32674 30046 32676 30098
rect 32172 29988 32228 29998
rect 32172 29894 32228 29932
rect 32396 29986 32452 29998
rect 32396 29934 32398 29986
rect 32450 29934 32452 29986
rect 32172 29316 32228 29326
rect 32172 29222 32228 29260
rect 32396 28532 32452 29934
rect 32620 28756 32676 30046
rect 33628 29426 33684 30156
rect 33628 29374 33630 29426
rect 33682 29374 33684 29426
rect 32732 29316 32788 29326
rect 32732 29222 32788 29260
rect 32620 28690 32676 28700
rect 32844 29202 32900 29214
rect 32844 29150 32846 29202
rect 32898 29150 32900 29202
rect 32844 28644 32900 29150
rect 33292 28868 33348 28878
rect 33292 28754 33348 28812
rect 33628 28868 33684 29374
rect 33628 28802 33684 28812
rect 33740 29314 33796 29326
rect 33740 29262 33742 29314
rect 33794 29262 33796 29314
rect 33292 28702 33294 28754
rect 33346 28702 33348 28754
rect 33292 28690 33348 28702
rect 33740 28756 33796 29262
rect 32844 28578 32900 28588
rect 32396 28196 32452 28476
rect 32396 28140 32676 28196
rect 32620 26962 32676 28140
rect 32620 26910 32622 26962
rect 32674 26910 32676 26962
rect 32732 27748 32788 27758
rect 32732 27076 32788 27692
rect 32732 26944 32788 27020
rect 33292 27188 33348 27198
rect 33292 27074 33348 27132
rect 33292 27022 33294 27074
rect 33346 27022 33348 27074
rect 33292 27010 33348 27022
rect 33740 27074 33796 28700
rect 33964 29204 34020 29214
rect 34188 29204 34244 29214
rect 33964 29202 34244 29204
rect 33964 29150 33966 29202
rect 34018 29150 34190 29202
rect 34242 29150 34244 29202
rect 33964 29148 34244 29150
rect 33964 27300 34020 29148
rect 34188 29138 34244 29148
rect 34188 28866 34244 28878
rect 34188 28814 34190 28866
rect 34242 28814 34244 28866
rect 34188 28754 34244 28814
rect 34188 28702 34190 28754
rect 34242 28702 34244 28754
rect 34188 28690 34244 28702
rect 33964 27234 34020 27244
rect 34076 28308 34132 28318
rect 34076 27298 34132 28252
rect 34076 27246 34078 27298
rect 34130 27246 34132 27298
rect 34076 27234 34132 27246
rect 33740 27022 33742 27074
rect 33794 27022 33796 27074
rect 33740 27010 33796 27022
rect 32620 26852 32676 26910
rect 34300 26908 34356 31388
rect 34636 29764 34692 33068
rect 34748 32788 34804 32798
rect 34972 32788 35028 33518
rect 35084 34130 35140 34142
rect 35084 34078 35086 34130
rect 35138 34078 35140 34130
rect 35084 33572 35140 34078
rect 35644 34018 35700 34030
rect 35644 33966 35646 34018
rect 35698 33966 35700 34018
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 33572 35252 33582
rect 35084 33570 35252 33572
rect 35084 33518 35198 33570
rect 35250 33518 35252 33570
rect 35084 33516 35252 33518
rect 34748 32786 35028 32788
rect 34748 32734 34750 32786
rect 34802 32734 35028 32786
rect 34748 32732 35028 32734
rect 35196 32788 35252 33516
rect 35420 33348 35476 33358
rect 35420 33254 35476 33292
rect 35644 33348 35700 33966
rect 35644 33282 35700 33292
rect 34748 32722 34804 32732
rect 35196 32722 35252 32732
rect 35532 33124 35588 33134
rect 35532 32786 35588 33068
rect 35532 32734 35534 32786
rect 35586 32734 35588 32786
rect 35532 32722 35588 32734
rect 35308 32674 35364 32686
rect 35308 32622 35310 32674
rect 35362 32622 35364 32674
rect 35196 32562 35252 32574
rect 35196 32510 35198 32562
rect 35250 32510 35252 32562
rect 35196 32452 35252 32510
rect 35308 32564 35364 32622
rect 35756 32564 35812 35532
rect 35868 35364 35924 35756
rect 35868 35298 35924 35308
rect 36092 35140 36148 38668
rect 36204 38668 36260 39116
rect 36316 39394 36372 39406
rect 36316 39342 36318 39394
rect 36370 39342 36372 39394
rect 36316 38948 36372 39342
rect 36540 39396 36596 40348
rect 36652 40292 36708 40302
rect 36652 40198 36708 40236
rect 36428 39060 36484 39070
rect 36540 39060 36596 39340
rect 36428 39058 36596 39060
rect 36428 39006 36430 39058
rect 36482 39006 36596 39058
rect 36428 39004 36596 39006
rect 36652 39394 36708 39406
rect 36652 39342 36654 39394
rect 36706 39342 36708 39394
rect 36428 38994 36484 39004
rect 36316 38882 36372 38892
rect 36204 38612 36484 38668
rect 35868 35084 36148 35140
rect 36204 37492 36260 37502
rect 35868 34356 35924 35084
rect 36204 35028 36260 37436
rect 36316 35586 36372 35598
rect 36316 35534 36318 35586
rect 36370 35534 36372 35586
rect 36316 35364 36372 35534
rect 36316 35298 36372 35308
rect 35868 34290 35924 34300
rect 35980 34972 36260 35028
rect 36316 35140 36372 35150
rect 35308 32508 35812 32564
rect 35196 32386 35252 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35756 31890 35812 32508
rect 35868 32452 35924 32462
rect 35868 32358 35924 32396
rect 35756 31838 35758 31890
rect 35810 31838 35812 31890
rect 35756 31826 35812 31838
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34412 29708 34692 29764
rect 34412 29650 34468 29708
rect 34412 29598 34414 29650
rect 34466 29598 34468 29650
rect 34412 29202 34468 29598
rect 34412 29150 34414 29202
rect 34466 29150 34468 29202
rect 34412 29138 34468 29150
rect 34524 29316 34580 29326
rect 34524 28866 34580 29260
rect 35756 29316 35812 29326
rect 35196 29036 35460 29046
rect 34524 28814 34526 28866
rect 34578 28814 34580 28866
rect 34524 28802 34580 28814
rect 34636 28980 34692 28990
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35756 28980 35812 29260
rect 34636 28756 34692 28924
rect 34636 28624 34692 28700
rect 35308 28868 35364 28878
rect 35308 28644 35364 28812
rect 35308 28530 35364 28588
rect 35308 28478 35310 28530
rect 35362 28478 35364 28530
rect 35308 28466 35364 28478
rect 35532 28756 35588 28766
rect 35532 28530 35588 28700
rect 35756 28754 35812 28924
rect 35980 28868 36036 34972
rect 36092 34692 36148 34702
rect 36092 34598 36148 34636
rect 36092 34356 36148 34366
rect 36092 34262 36148 34300
rect 36204 33906 36260 33918
rect 36204 33854 36206 33906
rect 36258 33854 36260 33906
rect 36092 33346 36148 33358
rect 36092 33294 36094 33346
rect 36146 33294 36148 33346
rect 36092 33124 36148 33294
rect 36092 33058 36148 33068
rect 36204 31444 36260 33854
rect 36316 33458 36372 35084
rect 36316 33406 36318 33458
rect 36370 33406 36372 33458
rect 36316 33394 36372 33406
rect 36428 33460 36484 38612
rect 36652 38612 36708 39342
rect 36652 38546 36708 38556
rect 36652 37938 36708 37950
rect 36652 37886 36654 37938
rect 36706 37886 36708 37938
rect 36540 37826 36596 37838
rect 36540 37774 36542 37826
rect 36594 37774 36596 37826
rect 36540 36820 36596 37774
rect 36652 37492 36708 37886
rect 36652 37426 36708 37436
rect 36540 36764 36708 36820
rect 36540 36596 36596 36606
rect 36540 34354 36596 36540
rect 36652 35588 36708 36764
rect 36652 35522 36708 35532
rect 36540 34302 36542 34354
rect 36594 34302 36596 34354
rect 36540 34290 36596 34302
rect 36652 35364 36708 35374
rect 36428 33394 36484 33404
rect 36540 33234 36596 33246
rect 36540 33182 36542 33234
rect 36594 33182 36596 33234
rect 36204 31378 36260 31388
rect 36316 32452 36372 32462
rect 36540 32452 36596 33182
rect 36652 33236 36708 35308
rect 36764 34242 36820 43260
rect 37100 43204 37156 43372
rect 36988 43148 37156 43204
rect 36764 34190 36766 34242
rect 36818 34190 36820 34242
rect 36764 34178 36820 34190
rect 36876 41524 36932 41534
rect 36876 34916 36932 41468
rect 36764 34020 36820 34030
rect 36764 33346 36820 33964
rect 36764 33294 36766 33346
rect 36818 33294 36820 33346
rect 36764 33282 36820 33294
rect 36652 33170 36708 33180
rect 36316 32450 36596 32452
rect 36316 32398 36318 32450
rect 36370 32398 36596 32450
rect 36316 32396 36596 32398
rect 35980 28812 36148 28868
rect 35756 28702 35758 28754
rect 35810 28702 35812 28754
rect 35756 28690 35812 28702
rect 35532 28478 35534 28530
rect 35586 28478 35588 28530
rect 35532 28466 35588 28478
rect 35980 28642 36036 28654
rect 35980 28590 35982 28642
rect 36034 28590 36036 28642
rect 35420 28420 35476 28430
rect 35420 28326 35476 28364
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35980 26964 36036 28590
rect 36092 27748 36148 28812
rect 36316 28308 36372 32396
rect 36876 31948 36932 34860
rect 36988 34468 37044 43148
rect 37212 40404 37268 44942
rect 37660 43540 37716 45612
rect 37772 45666 37828 49756
rect 39004 48692 39060 50764
rect 39116 50754 39172 50764
rect 39452 50484 39508 50988
rect 39452 50390 39508 50428
rect 39004 48626 39060 48636
rect 37996 48242 38052 48254
rect 37996 48190 37998 48242
rect 38050 48190 38052 48242
rect 37996 48132 38052 48190
rect 37996 48066 38052 48076
rect 38556 48132 38612 48142
rect 38556 48038 38612 48076
rect 37772 45614 37774 45666
rect 37826 45614 37828 45666
rect 37772 45602 37828 45614
rect 37884 48018 37940 48030
rect 37884 47966 37886 48018
rect 37938 47966 37940 48018
rect 37884 45668 37940 47966
rect 38332 47124 38388 47134
rect 38332 46114 38388 47068
rect 38332 46062 38334 46114
rect 38386 46062 38388 46114
rect 38332 46050 38388 46062
rect 37884 45574 37940 45612
rect 37996 45892 38052 45902
rect 37772 44996 37828 45006
rect 37772 44902 37828 44940
rect 37660 43474 37716 43484
rect 37996 43428 38052 45836
rect 38556 45890 38612 45902
rect 38556 45838 38558 45890
rect 38610 45838 38612 45890
rect 38556 45332 38612 45838
rect 39004 45668 39060 45678
rect 39004 45574 39060 45612
rect 38556 45266 38612 45276
rect 38220 45220 38276 45230
rect 39564 45220 39620 52780
rect 39900 53506 39956 53518
rect 39900 53454 39902 53506
rect 39954 53454 39956 53506
rect 39900 52164 39956 53454
rect 40012 53508 40068 53518
rect 40012 53414 40068 53452
rect 40684 53508 40740 53518
rect 40684 53414 40740 53452
rect 40796 53396 40852 53406
rect 40796 52836 40852 53340
rect 39900 52098 39956 52108
rect 40684 52834 40852 52836
rect 40684 52782 40798 52834
rect 40850 52782 40852 52834
rect 40684 52780 40852 52782
rect 40124 51604 40180 51614
rect 39788 51602 40180 51604
rect 39788 51550 40126 51602
rect 40178 51550 40180 51602
rect 39788 51548 40180 51550
rect 39788 50818 39844 51548
rect 40124 51538 40180 51548
rect 40236 51492 40292 51502
rect 39900 51378 39956 51390
rect 39900 51326 39902 51378
rect 39954 51326 39956 51378
rect 39900 51268 39956 51326
rect 40236 51378 40292 51436
rect 40236 51326 40238 51378
rect 40290 51326 40292 51378
rect 39900 51202 39956 51212
rect 40012 51266 40068 51278
rect 40012 51214 40014 51266
rect 40066 51214 40068 51266
rect 39788 50766 39790 50818
rect 39842 50766 39844 50818
rect 39788 50754 39844 50766
rect 40012 50820 40068 51214
rect 40236 51044 40292 51326
rect 40684 51380 40740 52780
rect 40796 52770 40852 52780
rect 40684 51314 40740 51324
rect 40796 52164 40852 52174
rect 40796 51378 40852 52108
rect 41244 51604 41300 53676
rect 41580 53666 41636 53676
rect 41916 53730 41972 53742
rect 41916 53678 41918 53730
rect 41970 53678 41972 53730
rect 41468 53506 41524 53518
rect 41468 53454 41470 53506
rect 41522 53454 41524 53506
rect 41468 53396 41524 53454
rect 41692 53508 41748 53518
rect 41692 53414 41748 53452
rect 41468 53330 41524 53340
rect 41244 51538 41300 51548
rect 41468 52834 41524 52846
rect 41468 52782 41470 52834
rect 41522 52782 41524 52834
rect 41468 52612 41524 52782
rect 41916 52612 41972 53678
rect 42140 53730 42196 53742
rect 42140 53678 42142 53730
rect 42194 53678 42196 53730
rect 42140 53620 42196 53678
rect 42140 53554 42196 53564
rect 41468 52556 41972 52612
rect 41468 51492 41524 52556
rect 41468 51426 41524 51436
rect 40796 51326 40798 51378
rect 40850 51326 40852 51378
rect 40796 51314 40852 51326
rect 42476 51380 42532 51390
rect 41580 51266 41636 51278
rect 41580 51214 41582 51266
rect 41634 51214 41636 51266
rect 40572 51156 40628 51166
rect 41580 51156 41636 51214
rect 40572 51154 41636 51156
rect 40572 51102 40574 51154
rect 40626 51102 41636 51154
rect 40572 51100 41636 51102
rect 40572 51090 40628 51100
rect 40236 50978 40292 50988
rect 40012 50754 40068 50764
rect 40460 50820 40516 50830
rect 40460 50726 40516 50764
rect 40124 50706 40180 50718
rect 40124 50654 40126 50706
rect 40178 50654 40180 50706
rect 40124 47124 40180 50654
rect 40124 47058 40180 47068
rect 40236 50484 40292 50494
rect 40236 46900 40292 50428
rect 40908 50484 40964 50494
rect 40908 50390 40964 50428
rect 40124 46844 40292 46900
rect 39900 45332 39956 45342
rect 39900 45238 39956 45276
rect 39788 45220 39844 45230
rect 39564 45218 39844 45220
rect 39564 45166 39790 45218
rect 39842 45166 39844 45218
rect 39564 45164 39844 45166
rect 38220 45126 38276 45164
rect 39788 44548 39844 45164
rect 40012 44996 40068 45006
rect 40012 44902 40068 44940
rect 40012 44548 40068 44558
rect 39788 44546 40068 44548
rect 39788 44494 40014 44546
rect 40066 44494 40068 44546
rect 39788 44492 40068 44494
rect 40012 44482 40068 44492
rect 40124 43708 40180 46844
rect 41580 46452 41636 51100
rect 42140 51266 42196 51278
rect 42140 51214 42142 51266
rect 42194 51214 42196 51266
rect 42140 51156 42196 51214
rect 42140 51090 42196 51100
rect 42476 51266 42532 51324
rect 42476 51214 42478 51266
rect 42530 51214 42532 51266
rect 42476 48132 42532 51214
rect 42476 48066 42532 48076
rect 41580 46386 41636 46396
rect 41804 46676 41860 46686
rect 41804 46562 41860 46620
rect 41804 46510 41806 46562
rect 41858 46510 41860 46562
rect 41020 45780 41076 45790
rect 40348 45668 40404 45678
rect 40348 45666 40740 45668
rect 40348 45614 40350 45666
rect 40402 45614 40740 45666
rect 40348 45612 40740 45614
rect 40348 45602 40404 45612
rect 40684 45218 40740 45612
rect 40796 45444 40852 45454
rect 40796 45330 40852 45388
rect 40796 45278 40798 45330
rect 40850 45278 40852 45330
rect 40796 45266 40852 45278
rect 40684 45166 40686 45218
rect 40738 45166 40740 45218
rect 37996 43362 38052 43372
rect 39676 43652 40180 43708
rect 40236 44546 40292 44558
rect 40236 44494 40238 44546
rect 40290 44494 40292 44546
rect 40236 44098 40292 44494
rect 40236 44046 40238 44098
rect 40290 44046 40292 44098
rect 37324 43316 37380 43326
rect 37324 43222 37380 43260
rect 37548 43314 37604 43326
rect 37548 43262 37550 43314
rect 37602 43262 37604 43314
rect 37548 41636 37604 43262
rect 37548 41570 37604 41580
rect 37660 42868 37716 42878
rect 37660 41300 37716 42812
rect 37660 41234 37716 41244
rect 37884 41972 37940 41982
rect 37884 41298 37940 41916
rect 37884 41246 37886 41298
rect 37938 41246 37940 41298
rect 37548 40964 37604 40974
rect 37548 40870 37604 40908
rect 37884 40852 37940 41246
rect 39676 41748 39732 43652
rect 39228 41076 39284 41086
rect 37100 40348 37268 40404
rect 37548 40402 37604 40414
rect 37548 40350 37550 40402
rect 37602 40350 37604 40402
rect 37100 36372 37156 40348
rect 37212 40178 37268 40190
rect 37212 40126 37214 40178
rect 37266 40126 37268 40178
rect 37212 36596 37268 40126
rect 37548 40068 37604 40350
rect 37884 40402 37940 40796
rect 37884 40350 37886 40402
rect 37938 40350 37940 40402
rect 37884 40338 37940 40350
rect 38556 40964 38612 40974
rect 38556 40628 38612 40908
rect 38556 40402 38612 40572
rect 38556 40350 38558 40402
rect 38610 40350 38612 40402
rect 38556 40338 38612 40350
rect 38780 40852 38836 40862
rect 38780 40514 38836 40796
rect 38780 40462 38782 40514
rect 38834 40462 38836 40514
rect 38780 40404 38836 40462
rect 38780 40338 38836 40348
rect 37436 39732 37492 39742
rect 37548 39732 37604 40012
rect 38556 39844 38612 39854
rect 37436 39730 37604 39732
rect 37436 39678 37438 39730
rect 37490 39678 37604 39730
rect 37436 39676 37604 39678
rect 38332 39732 38388 39742
rect 37436 39666 37492 39676
rect 38332 39638 38388 39676
rect 38108 39620 38164 39630
rect 38108 39526 38164 39564
rect 38556 39618 38612 39788
rect 38556 39566 38558 39618
rect 38610 39566 38612 39618
rect 38556 39554 38612 39566
rect 38780 39508 38836 39518
rect 38780 39414 38836 39452
rect 39228 39508 39284 41020
rect 39228 39414 39284 39452
rect 39228 39058 39284 39070
rect 39228 39006 39230 39058
rect 39282 39006 39284 39058
rect 39116 38948 39172 38958
rect 39116 38854 39172 38892
rect 38556 38836 38612 38846
rect 39004 38836 39060 38846
rect 38556 38834 39060 38836
rect 38556 38782 38558 38834
rect 38610 38782 39006 38834
rect 39058 38782 39060 38834
rect 38556 38780 39060 38782
rect 38556 38724 38612 38780
rect 39004 38770 39060 38780
rect 38556 38658 38612 38668
rect 37212 36530 37268 36540
rect 38444 37940 38500 37950
rect 37100 36306 37156 36316
rect 37436 36372 37492 36382
rect 36988 34402 37044 34412
rect 37100 35812 37156 35822
rect 36988 34020 37044 34030
rect 36988 33926 37044 33964
rect 37100 32900 37156 35756
rect 37436 34354 37492 36316
rect 38220 35812 38276 35822
rect 38220 35718 38276 35756
rect 37436 34302 37438 34354
rect 37490 34302 37492 34354
rect 37436 33906 37492 34302
rect 38108 35476 38164 35486
rect 37884 34020 37940 34030
rect 37436 33854 37438 33906
rect 37490 33854 37492 33906
rect 37436 33842 37492 33854
rect 37660 34018 37940 34020
rect 37660 33966 37886 34018
rect 37938 33966 37940 34018
rect 37660 33964 37940 33966
rect 37100 32834 37156 32844
rect 37324 33236 37380 33246
rect 37212 32788 37268 32798
rect 37212 32694 37268 32732
rect 37324 32674 37380 33180
rect 37324 32622 37326 32674
rect 37378 32622 37380 32674
rect 37324 32610 37380 32622
rect 37660 33122 37716 33964
rect 37884 33954 37940 33964
rect 37996 33906 38052 33918
rect 37996 33854 37998 33906
rect 38050 33854 38052 33906
rect 37996 33346 38052 33854
rect 37996 33294 37998 33346
rect 38050 33294 38052 33346
rect 37996 33282 38052 33294
rect 37660 33070 37662 33122
rect 37714 33070 37716 33122
rect 36764 31892 36932 31948
rect 36988 32452 37044 32462
rect 36764 28980 36820 31892
rect 36876 31780 36932 31790
rect 36876 31686 36932 31724
rect 36988 30996 37044 32396
rect 36988 30930 37044 30940
rect 37436 30882 37492 30894
rect 37436 30830 37438 30882
rect 37490 30830 37492 30882
rect 37436 30212 37492 30830
rect 37436 30146 37492 30156
rect 36764 28914 36820 28924
rect 37660 28756 37716 33070
rect 37772 33122 37828 33134
rect 37772 33070 37774 33122
rect 37826 33070 37828 33122
rect 37772 31668 37828 33070
rect 37884 33122 37940 33134
rect 37884 33070 37886 33122
rect 37938 33070 37940 33122
rect 37884 32788 37940 33070
rect 37884 32722 37940 32732
rect 38108 32450 38164 35420
rect 38332 33572 38388 33582
rect 38332 33478 38388 33516
rect 38220 33012 38276 33022
rect 38220 32786 38276 32956
rect 38220 32734 38222 32786
rect 38274 32734 38276 32786
rect 38220 32722 38276 32734
rect 38444 32564 38500 37884
rect 39116 37940 39172 37950
rect 39116 37846 39172 37884
rect 38668 35588 38724 35598
rect 38668 35494 38724 35532
rect 39116 35252 39172 35262
rect 39116 34690 39172 35196
rect 39116 34638 39118 34690
rect 39170 34638 39172 34690
rect 39116 34468 39172 34638
rect 39116 34402 39172 34412
rect 39228 33908 39284 39006
rect 39452 38052 39508 38062
rect 39676 38052 39732 41692
rect 39900 41636 39956 41646
rect 39900 40290 39956 41580
rect 39900 40238 39902 40290
rect 39954 40238 39956 40290
rect 39900 40226 39956 40238
rect 40012 40964 40068 40974
rect 40012 40514 40068 40908
rect 40236 40964 40292 44046
rect 40236 40898 40292 40908
rect 40572 40964 40628 40974
rect 40012 40462 40014 40514
rect 40066 40462 40068 40514
rect 39900 39620 39956 39630
rect 39900 39526 39956 39564
rect 40012 38612 40068 40462
rect 40460 40740 40516 40750
rect 40236 40404 40292 40414
rect 40236 40290 40292 40348
rect 40236 40238 40238 40290
rect 40290 40238 40292 40290
rect 40236 40226 40292 40238
rect 40460 39618 40516 40684
rect 40572 40628 40628 40908
rect 40684 40852 40740 45166
rect 40684 40786 40740 40796
rect 40684 40628 40740 40638
rect 40572 40626 40740 40628
rect 40572 40574 40686 40626
rect 40738 40574 40740 40626
rect 40572 40572 40740 40574
rect 40684 40562 40740 40572
rect 40796 40180 40852 40190
rect 40684 40068 40740 40078
rect 40572 39844 40628 39854
rect 40572 39750 40628 39788
rect 40460 39566 40462 39618
rect 40514 39566 40516 39618
rect 40460 39554 40516 39566
rect 40572 39620 40628 39630
rect 40684 39620 40740 40012
rect 40628 39564 40740 39620
rect 40572 39506 40628 39564
rect 40572 39454 40574 39506
rect 40626 39454 40628 39506
rect 40572 39442 40628 39454
rect 40684 39396 40740 39406
rect 40572 38948 40628 38958
rect 40572 38854 40628 38892
rect 40684 38834 40740 39340
rect 40684 38782 40686 38834
rect 40738 38782 40740 38834
rect 40684 38770 40740 38782
rect 39900 38556 40068 38612
rect 39452 38050 39732 38052
rect 39452 37998 39454 38050
rect 39506 37998 39732 38050
rect 39452 37996 39732 37998
rect 39452 37986 39508 37996
rect 39452 37828 39508 37838
rect 39452 37734 39508 37772
rect 39676 37156 39732 37996
rect 39788 38052 39844 38062
rect 39788 37958 39844 37996
rect 39788 37156 39844 37166
rect 39676 37154 39844 37156
rect 39676 37102 39790 37154
rect 39842 37102 39844 37154
rect 39676 37100 39844 37102
rect 39788 36932 39844 37100
rect 39788 36866 39844 36876
rect 39564 36260 39620 36270
rect 39564 35812 39620 36204
rect 39676 36148 39732 36158
rect 39676 35922 39732 36092
rect 39676 35870 39678 35922
rect 39730 35870 39732 35922
rect 39676 35858 39732 35870
rect 39564 35718 39620 35756
rect 39788 35698 39844 35710
rect 39788 35646 39790 35698
rect 39842 35646 39844 35698
rect 39788 35588 39844 35646
rect 39788 35522 39844 35532
rect 39900 35364 39956 38556
rect 40236 37938 40292 37950
rect 40236 37886 40238 37938
rect 40290 37886 40292 37938
rect 40236 37828 40292 37886
rect 40236 37772 40740 37828
rect 40460 37378 40516 37390
rect 40460 37326 40462 37378
rect 40514 37326 40516 37378
rect 40460 37268 40516 37326
rect 40684 37378 40740 37772
rect 40684 37326 40686 37378
rect 40738 37326 40740 37378
rect 40684 37314 40740 37326
rect 40124 36484 40180 36494
rect 40012 36372 40068 36382
rect 40012 36278 40068 36316
rect 40012 35588 40068 35598
rect 40012 35494 40068 35532
rect 39900 35308 40068 35364
rect 40012 34804 40068 35308
rect 40124 34916 40180 36428
rect 40460 35700 40516 37212
rect 40572 37154 40628 37166
rect 40572 37102 40574 37154
rect 40626 37102 40628 37154
rect 40572 36708 40628 37102
rect 40572 36642 40628 36652
rect 40796 36594 40852 40124
rect 40796 36542 40798 36594
rect 40850 36542 40852 36594
rect 40796 36530 40852 36542
rect 40908 38724 40964 38734
rect 40908 38050 40964 38668
rect 40908 37998 40910 38050
rect 40962 37998 40964 38050
rect 40684 36260 40740 36270
rect 40684 36166 40740 36204
rect 40908 36258 40964 37998
rect 40908 36206 40910 36258
rect 40962 36206 40964 36258
rect 40460 35644 40628 35700
rect 40236 35474 40292 35486
rect 40460 35476 40516 35486
rect 40236 35422 40238 35474
rect 40290 35422 40292 35474
rect 40236 35140 40292 35422
rect 40236 35074 40292 35084
rect 40348 35474 40516 35476
rect 40348 35422 40462 35474
rect 40514 35422 40516 35474
rect 40348 35420 40516 35422
rect 40236 34916 40292 34926
rect 40124 34914 40292 34916
rect 40124 34862 40238 34914
rect 40290 34862 40292 34914
rect 40124 34860 40292 34862
rect 40236 34850 40292 34860
rect 40012 34748 40180 34804
rect 39900 34690 39956 34702
rect 39900 34638 39902 34690
rect 39954 34638 39956 34690
rect 39900 34244 39956 34638
rect 39900 34178 39956 34188
rect 39228 33842 39284 33852
rect 40012 33458 40068 33470
rect 40012 33406 40014 33458
rect 40066 33406 40068 33458
rect 38108 32398 38110 32450
rect 38162 32398 38164 32450
rect 38108 32386 38164 32398
rect 38332 32508 38500 32564
rect 38556 33346 38612 33358
rect 38556 33294 38558 33346
rect 38610 33294 38612 33346
rect 38108 31780 38164 31790
rect 38332 31780 38388 32508
rect 38444 32340 38500 32350
rect 38444 32246 38500 32284
rect 38556 31948 38612 33294
rect 38892 33236 38948 33246
rect 38892 32786 38948 33180
rect 38892 32734 38894 32786
rect 38946 32734 38948 32786
rect 38892 32722 38948 32734
rect 39004 33122 39060 33134
rect 39004 33070 39006 33122
rect 39058 33070 39060 33122
rect 39004 33012 39060 33070
rect 39004 32116 39060 32956
rect 38556 31892 38724 31948
rect 38668 31826 38724 31836
rect 38556 31780 38612 31790
rect 38332 31778 38612 31780
rect 38332 31726 38558 31778
rect 38610 31726 38612 31778
rect 38332 31724 38612 31726
rect 39004 31780 39060 32060
rect 39564 33122 39620 33134
rect 39564 33070 39566 33122
rect 39618 33070 39620 33122
rect 39564 32786 39620 33070
rect 39564 32734 39566 32786
rect 39618 32734 39620 32786
rect 39228 31892 39284 31902
rect 39228 31798 39284 31836
rect 39116 31780 39172 31790
rect 39004 31778 39172 31780
rect 39004 31726 39118 31778
rect 39170 31726 39172 31778
rect 39004 31724 39172 31726
rect 38108 31686 38164 31724
rect 38556 31714 38612 31724
rect 39116 31714 39172 31724
rect 37772 31602 37828 31612
rect 37884 31666 37940 31678
rect 37884 31614 37886 31666
rect 37938 31614 37940 31666
rect 37884 31556 37940 31614
rect 37884 31490 37940 31500
rect 37996 31666 38052 31678
rect 37996 31614 37998 31666
rect 38050 31614 38052 31666
rect 37996 30212 38052 31614
rect 39452 31668 39508 31678
rect 39452 31574 39508 31612
rect 39564 31556 39620 32734
rect 39900 32676 39956 32686
rect 39900 32116 39956 32620
rect 40012 32228 40068 33406
rect 40124 32452 40180 34748
rect 40124 32358 40180 32396
rect 40012 32172 40180 32228
rect 39900 31890 39956 32060
rect 39900 31838 39902 31890
rect 39954 31838 39956 31890
rect 39900 31826 39956 31838
rect 40012 32004 40068 32014
rect 39564 31490 39620 31500
rect 39900 31444 39956 31454
rect 39900 31218 39956 31388
rect 39900 31166 39902 31218
rect 39954 31166 39956 31218
rect 39900 31154 39956 31166
rect 40012 31218 40068 31948
rect 40124 31444 40180 32172
rect 40348 32004 40404 35420
rect 40460 35410 40516 35420
rect 40572 35252 40628 35644
rect 40348 31938 40404 31948
rect 40460 34914 40516 34926
rect 40460 34862 40462 34914
rect 40514 34862 40516 34914
rect 40124 31378 40180 31388
rect 40348 31668 40404 31678
rect 40348 31554 40404 31612
rect 40348 31502 40350 31554
rect 40402 31502 40404 31554
rect 40012 31166 40014 31218
rect 40066 31166 40068 31218
rect 40012 31154 40068 31166
rect 40124 30884 40180 30894
rect 40124 30790 40180 30828
rect 37996 30146 38052 30156
rect 37660 28690 37716 28700
rect 38108 29204 38164 29214
rect 38108 28644 38164 29148
rect 39340 28868 39396 28878
rect 38108 28550 38164 28588
rect 38556 28642 38612 28654
rect 38556 28590 38558 28642
rect 38610 28590 38612 28642
rect 36316 28242 36372 28252
rect 38556 28308 38612 28590
rect 38556 28242 38612 28252
rect 39116 28530 39172 28542
rect 39116 28478 39118 28530
rect 39170 28478 39172 28530
rect 39116 28308 39172 28478
rect 39340 28530 39396 28812
rect 39564 28644 39620 28654
rect 39564 28550 39620 28588
rect 39900 28644 39956 28682
rect 39900 28578 39956 28588
rect 39340 28478 39342 28530
rect 39394 28478 39396 28530
rect 39340 28466 39396 28478
rect 39116 28242 39172 28252
rect 39900 28418 39956 28430
rect 39900 28366 39902 28418
rect 39954 28366 39956 28418
rect 36092 27682 36148 27692
rect 34300 26852 35140 26908
rect 35980 26898 36036 26908
rect 32172 26796 32676 26852
rect 32172 26514 32228 26796
rect 32172 26462 32174 26514
rect 32226 26462 32228 26514
rect 32172 26450 32228 26462
rect 31612 8372 31892 8428
rect 32508 24052 32564 24062
rect 29372 3444 29428 3454
rect 29820 3444 29876 3454
rect 29372 3442 29876 3444
rect 29372 3390 29374 3442
rect 29426 3390 29822 3442
rect 29874 3390 29876 3442
rect 29372 3388 29876 3390
rect 29372 3378 29428 3388
rect 28140 3266 28196 3276
rect 20748 728 21000 800
rect 20776 200 21000 728
rect 23464 200 23688 800
rect 26824 728 27076 800
rect 29484 800 29540 3388
rect 29820 3378 29876 3388
rect 30156 3332 30212 3342
rect 30156 3238 30212 3276
rect 31612 3332 31668 8372
rect 32508 3666 32564 23996
rect 35084 8428 35140 26852
rect 39900 26404 39956 28366
rect 39900 26338 39956 26348
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 32508 3614 32510 3666
rect 32562 3614 32564 3666
rect 32508 3556 32564 3614
rect 34748 8372 35140 8428
rect 34748 4562 34804 8372
rect 40348 8148 40404 31502
rect 40460 31556 40516 34862
rect 40572 34132 40628 35196
rect 40572 34066 40628 34076
rect 40908 33348 40964 36206
rect 40908 33282 40964 33292
rect 40460 31490 40516 31500
rect 40684 32450 40740 32462
rect 40684 32398 40686 32450
rect 40738 32398 40740 32450
rect 40684 32340 40740 32398
rect 40572 31444 40628 31454
rect 40572 31218 40628 31388
rect 40572 31166 40574 31218
rect 40626 31166 40628 31218
rect 40572 31154 40628 31166
rect 40460 28644 40516 28654
rect 40460 28550 40516 28588
rect 40348 8082 40404 8092
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34748 4510 34750 4562
rect 34802 4510 34804 4562
rect 33180 3556 33236 3566
rect 32508 3554 33236 3556
rect 32508 3502 33182 3554
rect 33234 3502 33236 3554
rect 32508 3500 33236 3502
rect 34748 3556 34804 4510
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35756 3666 35812 3678
rect 35756 3614 35758 3666
rect 35810 3614 35812 3666
rect 35084 3556 35140 3566
rect 34748 3554 35140 3556
rect 34748 3502 35086 3554
rect 35138 3502 35140 3554
rect 34748 3500 35140 3502
rect 33180 3490 33236 3500
rect 35084 3490 35140 3500
rect 31612 3266 31668 3276
rect 32396 3444 32452 3454
rect 32396 800 32452 3388
rect 34076 3444 34132 3454
rect 34076 3350 34132 3388
rect 35756 800 35812 3614
rect 40684 3220 40740 32284
rect 41020 30324 41076 45724
rect 41244 44996 41300 45006
rect 41132 40740 41188 40750
rect 41132 39730 41188 40684
rect 41132 39678 41134 39730
rect 41186 39678 41188 39730
rect 41132 39666 41188 39678
rect 41132 38164 41188 38174
rect 41132 37156 41188 38108
rect 41132 37090 41188 37100
rect 41132 36484 41188 36494
rect 41132 36390 41188 36428
rect 41244 31948 41300 44940
rect 41580 44996 41636 45006
rect 41580 44902 41636 44940
rect 41804 41972 41860 46510
rect 42364 46564 42420 46574
rect 42364 46470 42420 46508
rect 41804 41906 41860 41916
rect 41916 45444 41972 45454
rect 41804 41074 41860 41086
rect 41804 41022 41806 41074
rect 41858 41022 41860 41074
rect 41468 40404 41524 40414
rect 41468 40310 41524 40348
rect 41804 39844 41860 41022
rect 41916 41074 41972 45388
rect 42588 43708 42644 56028
rect 42812 53620 42868 53630
rect 42812 53526 42868 53564
rect 42700 53060 42756 53070
rect 42700 52966 42756 53004
rect 43372 53060 43428 53070
rect 43260 52724 43316 52734
rect 42812 52722 43316 52724
rect 42812 52670 43262 52722
rect 43314 52670 43316 52722
rect 42812 52668 43316 52670
rect 42588 43652 42756 43708
rect 42140 41188 42196 41198
rect 42588 41188 42644 41198
rect 42140 41186 42644 41188
rect 42140 41134 42142 41186
rect 42194 41134 42590 41186
rect 42642 41134 42644 41186
rect 42140 41132 42644 41134
rect 42140 41122 42196 41132
rect 42588 41122 42644 41132
rect 41916 41022 41918 41074
rect 41970 41022 41972 41074
rect 41916 41010 41972 41022
rect 42700 40964 42756 43652
rect 42812 42532 42868 52668
rect 43260 52658 43316 52668
rect 43148 51378 43204 51390
rect 43148 51326 43150 51378
rect 43202 51326 43204 51378
rect 43036 51266 43092 51278
rect 43036 51214 43038 51266
rect 43090 51214 43092 51266
rect 43036 50820 43092 51214
rect 43148 51156 43204 51326
rect 43148 51090 43204 51100
rect 43036 50754 43092 50764
rect 43372 50036 43428 53004
rect 43596 52836 43652 52846
rect 43596 52742 43652 52780
rect 44044 52836 44100 52846
rect 44044 52742 44100 52780
rect 43484 51380 43540 51390
rect 43484 51286 43540 51324
rect 43596 50036 43652 50046
rect 43260 49980 43596 50036
rect 43036 48020 43092 48030
rect 43036 46898 43092 47964
rect 43036 46846 43038 46898
rect 43090 46846 43092 46898
rect 43036 46834 43092 46846
rect 42924 46676 42980 46686
rect 42924 46582 42980 46620
rect 43148 46674 43204 46686
rect 43148 46622 43150 46674
rect 43202 46622 43204 46674
rect 43148 45444 43204 46622
rect 43148 45378 43204 45388
rect 42812 42476 43092 42532
rect 42812 41300 42868 41310
rect 42812 41206 42868 41244
rect 42476 40908 42756 40964
rect 42924 41186 42980 41198
rect 42924 41134 42926 41186
rect 42978 41134 42980 41186
rect 41804 39778 41860 39788
rect 42028 40852 42084 40862
rect 42028 39730 42084 40796
rect 42028 39678 42030 39730
rect 42082 39678 42084 39730
rect 42028 39666 42084 39678
rect 42140 40740 42196 40750
rect 42140 40402 42196 40684
rect 42140 40350 42142 40402
rect 42194 40350 42196 40402
rect 42140 39732 42196 40350
rect 42476 40626 42532 40908
rect 42476 40574 42478 40626
rect 42530 40574 42532 40626
rect 42476 40292 42532 40574
rect 42700 40740 42756 40750
rect 42700 40626 42756 40684
rect 42700 40574 42702 40626
rect 42754 40574 42756 40626
rect 42700 40562 42756 40574
rect 42476 40226 42532 40236
rect 42812 40180 42868 40190
rect 42924 40180 42980 41134
rect 42812 40178 42980 40180
rect 42812 40126 42814 40178
rect 42866 40126 42980 40178
rect 42812 40124 42980 40126
rect 42476 39732 42532 39742
rect 42140 39730 42532 39732
rect 42140 39678 42478 39730
rect 42530 39678 42532 39730
rect 42140 39676 42532 39678
rect 42476 39666 42532 39676
rect 42812 39620 42868 40124
rect 42812 39554 42868 39564
rect 41580 39396 41636 39406
rect 41580 39302 41636 39340
rect 41916 38948 41972 38958
rect 41580 38724 41636 38734
rect 41580 38630 41636 38668
rect 41916 38722 41972 38892
rect 41916 38670 41918 38722
rect 41970 38670 41972 38722
rect 41692 38164 41748 38174
rect 41692 38070 41748 38108
rect 41468 37268 41524 37278
rect 41468 37174 41524 37212
rect 41692 36932 41748 36942
rect 41356 36708 41412 36718
rect 41356 36614 41412 36652
rect 41580 36596 41636 36606
rect 41580 36502 41636 36540
rect 41692 35364 41748 36876
rect 41916 36932 41972 38670
rect 42140 38052 42196 38062
rect 42140 37958 42196 37996
rect 41916 36866 41972 36876
rect 42476 37492 42532 37502
rect 42476 36706 42532 37436
rect 43036 36820 43092 42476
rect 43260 41300 43316 49980
rect 43596 49904 43652 49980
rect 44268 50036 44324 50046
rect 44940 50036 44996 56140
rect 46620 56194 46676 56206
rect 46620 56142 46622 56194
rect 46674 56142 46676 56194
rect 46620 55468 46676 56142
rect 46844 56082 46900 56364
rect 46844 56030 46846 56082
rect 46898 56030 46900 56082
rect 46844 56018 46900 56030
rect 49532 56084 49588 56094
rect 49532 55990 49588 56028
rect 49868 55972 49924 59200
rect 52332 59200 52584 59304
rect 55720 59304 55944 59800
rect 55720 59200 55972 59304
rect 52332 56642 52388 59200
rect 52332 56590 52334 56642
rect 52386 56590 52388 56642
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 52108 56308 52164 56318
rect 52332 56308 52388 56590
rect 52108 56306 52388 56308
rect 52108 56254 52110 56306
rect 52162 56254 52388 56306
rect 52108 56252 52388 56254
rect 53004 56642 53060 56654
rect 53004 56590 53006 56642
rect 53058 56590 53060 56642
rect 52108 56242 52164 56252
rect 52780 56196 52836 56206
rect 52780 56102 52836 56140
rect 49980 56084 50036 56094
rect 49980 55990 50036 56028
rect 53004 56082 53060 56590
rect 55132 56308 55188 56318
rect 55132 56214 55188 56252
rect 55916 56308 55972 59200
rect 53004 56030 53006 56082
rect 53058 56030 53060 56082
rect 53004 56018 53060 56030
rect 55580 56194 55636 56206
rect 55580 56142 55582 56194
rect 55634 56142 55636 56194
rect 49868 55906 49924 55916
rect 50652 55972 50708 55982
rect 50652 55878 50708 55916
rect 46508 55412 46676 55468
rect 45612 53618 45668 53630
rect 45612 53566 45614 53618
rect 45666 53566 45668 53618
rect 45500 53508 45556 53518
rect 45612 53508 45668 53566
rect 46060 53508 46116 53518
rect 45612 53506 46116 53508
rect 45612 53454 46062 53506
rect 46114 53454 46116 53506
rect 45612 53452 46116 53454
rect 45500 53414 45556 53452
rect 46060 52276 46116 53452
rect 46060 50708 46116 52220
rect 46060 50642 46116 50652
rect 44268 49942 44324 49980
rect 44492 50034 44996 50036
rect 44492 49982 44942 50034
rect 44994 49982 44996 50034
rect 44492 49980 44996 49982
rect 44492 49922 44548 49980
rect 44940 49970 44996 49980
rect 44492 49870 44494 49922
rect 44546 49870 44548 49922
rect 44492 49858 44548 49870
rect 44156 49588 44212 49598
rect 43820 49586 44212 49588
rect 43820 49534 44158 49586
rect 44210 49534 44212 49586
rect 43820 49532 44212 49534
rect 43820 46674 43876 49532
rect 44156 49522 44212 49532
rect 43820 46622 43822 46674
rect 43874 46622 43876 46674
rect 43820 46610 43876 46622
rect 43148 41244 43316 41300
rect 43372 46564 43428 46574
rect 43148 40628 43204 41244
rect 43260 41076 43316 41086
rect 43260 40982 43316 41020
rect 43148 40572 43316 40628
rect 43148 40402 43204 40414
rect 43148 40350 43150 40402
rect 43202 40350 43204 40402
rect 43148 40292 43204 40350
rect 43148 40226 43204 40236
rect 43036 36754 43092 36764
rect 43260 36708 43316 40572
rect 43372 40516 43428 46508
rect 43596 46450 43652 46462
rect 43596 46398 43598 46450
rect 43650 46398 43652 46450
rect 43596 41300 43652 46398
rect 46508 45220 46564 55412
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 51436 53620 51492 53630
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 51436 52386 51492 53564
rect 55580 52836 55636 56142
rect 55916 56194 55972 56252
rect 55916 56142 55918 56194
rect 55970 56142 55972 56194
rect 55916 56130 55972 56142
rect 57708 59276 58324 59332
rect 58408 59304 58632 59800
rect 57708 56194 57764 59276
rect 58268 59220 58324 59276
rect 58380 59220 58632 59304
rect 58268 59200 58632 59220
rect 58268 59164 58436 59200
rect 57708 56142 57710 56194
rect 57762 56142 57764 56194
rect 57708 56130 57764 56142
rect 57820 57764 57876 57774
rect 56812 56084 56868 56094
rect 56588 56082 56868 56084
rect 56588 56030 56814 56082
rect 56866 56030 56868 56082
rect 56588 56028 56868 56030
rect 55580 52770 55636 52780
rect 55804 55522 55860 55534
rect 55804 55470 55806 55522
rect 55858 55470 55860 55522
rect 55804 55074 55860 55470
rect 56588 55522 56644 56028
rect 56812 56018 56868 56028
rect 56588 55470 56590 55522
rect 56642 55470 56644 55522
rect 56588 55458 56644 55470
rect 57820 55410 57876 57708
rect 57820 55358 57822 55410
rect 57874 55358 57876 55410
rect 57820 55346 57876 55358
rect 58044 55412 58100 55422
rect 56812 55300 56868 55310
rect 55804 55022 55806 55074
rect 55858 55022 55860 55074
rect 51436 52334 51438 52386
rect 51490 52334 51492 52386
rect 51436 52322 51492 52334
rect 52668 52276 52724 52286
rect 52668 52182 52724 52220
rect 51772 52164 51828 52174
rect 51772 52070 51828 52108
rect 52220 52162 52276 52174
rect 52220 52110 52222 52162
rect 52274 52110 52276 52162
rect 51548 51940 51604 51950
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 47068 50708 47124 50718
rect 46620 48580 46676 48590
rect 46620 48466 46676 48524
rect 46620 48414 46622 48466
rect 46674 48414 46676 48466
rect 46620 47572 46676 48414
rect 47068 48466 47124 50652
rect 51548 50596 51604 51884
rect 52220 51940 52276 52110
rect 53452 52164 53508 52174
rect 53452 52070 53508 52108
rect 53564 52162 53620 52174
rect 53564 52110 53566 52162
rect 53618 52110 53620 52162
rect 52220 51874 52276 51884
rect 53564 51716 53620 52110
rect 54124 52164 54180 52174
rect 54124 52070 54180 52108
rect 51548 50530 51604 50540
rect 53116 51660 53620 51716
rect 53116 51602 53172 51660
rect 53116 51550 53118 51602
rect 53170 51550 53172 51602
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 47068 48414 47070 48466
rect 47122 48414 47124 48466
rect 47068 48356 47124 48414
rect 46844 47572 46900 47582
rect 46620 47570 46900 47572
rect 46620 47518 46846 47570
rect 46898 47518 46900 47570
rect 46620 47516 46900 47518
rect 47068 47572 47124 48300
rect 47516 48802 47572 48814
rect 47516 48750 47518 48802
rect 47570 48750 47572 48802
rect 47516 48692 47572 48750
rect 49084 48804 49140 48814
rect 47516 48244 47572 48636
rect 48188 48692 48244 48702
rect 47516 48178 47572 48188
rect 47852 48580 47908 48590
rect 47852 48244 47908 48524
rect 48076 48356 48132 48366
rect 47852 48242 48020 48244
rect 47852 48190 47854 48242
rect 47906 48190 48020 48242
rect 47852 48188 48020 48190
rect 47852 48178 47908 48188
rect 47292 47572 47348 47582
rect 47068 47570 47348 47572
rect 47068 47518 47294 47570
rect 47346 47518 47348 47570
rect 47068 47516 47348 47518
rect 46844 47506 46900 47516
rect 47292 47506 47348 47516
rect 47964 47460 48020 48188
rect 48076 48132 48132 48300
rect 48188 48354 48244 48636
rect 48188 48302 48190 48354
rect 48242 48302 48244 48354
rect 48188 48290 48244 48302
rect 48076 48076 48356 48132
rect 48076 47460 48132 47470
rect 47964 47458 48132 47460
rect 47964 47406 48078 47458
rect 48130 47406 48132 47458
rect 47964 47404 48132 47406
rect 48076 47394 48132 47404
rect 48300 47458 48356 48076
rect 48636 48020 48692 48030
rect 48300 47406 48302 47458
rect 48354 47406 48356 47458
rect 48300 47394 48356 47406
rect 48524 48018 48692 48020
rect 48524 47966 48638 48018
rect 48690 47966 48692 48018
rect 48524 47964 48692 47966
rect 48412 47234 48468 47246
rect 48412 47182 48414 47234
rect 48466 47182 48468 47234
rect 48412 46788 48468 47182
rect 47964 46732 48468 46788
rect 47964 46674 48020 46732
rect 48524 46676 48580 47964
rect 48636 47954 48692 47964
rect 49084 47572 49140 48748
rect 53116 48804 53172 51550
rect 55804 51380 55860 55022
rect 56252 55298 56868 55300
rect 56252 55246 56814 55298
rect 56866 55246 56868 55298
rect 56252 55244 56868 55246
rect 56252 55074 56308 55244
rect 56812 55234 56868 55244
rect 56252 55022 56254 55074
rect 56306 55022 56308 55074
rect 56252 52164 56308 55022
rect 58044 54738 58100 55356
rect 58044 54686 58046 54738
rect 58098 54686 58100 54738
rect 58044 54674 58100 54686
rect 56252 52098 56308 52108
rect 55804 51314 55860 51324
rect 57260 50484 57316 50494
rect 57260 50390 57316 50428
rect 58044 50484 58100 50494
rect 58044 50390 58100 50428
rect 57708 50372 57764 50382
rect 53116 48738 53172 48748
rect 57596 50370 57764 50372
rect 57596 50318 57710 50370
rect 57762 50318 57764 50370
rect 57596 50316 57764 50318
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 48748 47570 49140 47572
rect 48748 47518 49086 47570
rect 49138 47518 49140 47570
rect 48748 47516 49140 47518
rect 48748 47458 48804 47516
rect 49084 47506 49140 47516
rect 48748 47406 48750 47458
rect 48802 47406 48804 47458
rect 48748 47394 48804 47406
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 47964 46622 47966 46674
rect 48018 46622 48020 46674
rect 47964 46610 48020 46622
rect 48076 46620 48580 46676
rect 47740 46564 47796 46574
rect 47740 46470 47796 46508
rect 48076 46562 48132 46620
rect 48076 46510 48078 46562
rect 48130 46510 48132 46562
rect 48076 46498 48132 46510
rect 48748 46564 48804 46574
rect 48748 46470 48804 46508
rect 50092 46564 50148 46574
rect 47628 46452 47684 46462
rect 47628 46358 47684 46396
rect 46508 45154 46564 45164
rect 45612 42642 45668 42654
rect 45612 42590 45614 42642
rect 45666 42590 45668 42642
rect 45500 42530 45556 42542
rect 45500 42478 45502 42530
rect 45554 42478 45556 42530
rect 43596 41234 43652 41244
rect 44156 41972 44212 41982
rect 43820 40964 43876 40974
rect 43820 40870 43876 40908
rect 43428 40460 43764 40516
rect 43372 40384 43428 40460
rect 43708 38724 43764 40460
rect 44156 39060 44212 41916
rect 45500 39396 45556 42478
rect 45276 39060 45332 39070
rect 44156 39058 45332 39060
rect 44156 39006 44158 39058
rect 44210 39006 45278 39058
rect 45330 39006 45332 39058
rect 44156 39004 45332 39006
rect 44156 38994 44212 39004
rect 42476 36654 42478 36706
rect 42530 36654 42532 36706
rect 42476 36642 42532 36654
rect 43148 36652 43316 36708
rect 43484 37492 43540 37502
rect 42140 36596 42196 36606
rect 42924 36596 42980 36606
rect 43148 36596 43204 36652
rect 42140 36502 42196 36540
rect 42588 36594 43204 36596
rect 42588 36542 42926 36594
rect 42978 36542 43204 36594
rect 42588 36540 43204 36542
rect 42252 36372 42308 36382
rect 42588 36372 42644 36540
rect 42924 36530 42980 36540
rect 42252 36370 42644 36372
rect 42252 36318 42254 36370
rect 42306 36318 42644 36370
rect 42252 36316 42644 36318
rect 42252 36306 42308 36316
rect 41804 35588 41860 35598
rect 41804 35586 41972 35588
rect 41804 35534 41806 35586
rect 41858 35534 41972 35586
rect 41804 35532 41972 35534
rect 41804 35522 41860 35532
rect 41804 35364 41860 35374
rect 41692 35308 41804 35364
rect 41020 30258 41076 30268
rect 41132 31892 41300 31948
rect 41692 33124 41748 33134
rect 41132 17556 41188 31892
rect 41692 31780 41748 33068
rect 41804 31948 41860 35308
rect 41916 33348 41972 35532
rect 42700 35028 42756 35038
rect 42028 33460 42084 33470
rect 42028 33366 42084 33404
rect 42476 33460 42532 33470
rect 41916 33254 41972 33292
rect 42140 32562 42196 32574
rect 42140 32510 42142 32562
rect 42194 32510 42196 32562
rect 41804 31892 41972 31948
rect 41804 31780 41860 31790
rect 41244 31778 41860 31780
rect 41244 31726 41806 31778
rect 41858 31726 41860 31778
rect 41244 31724 41860 31726
rect 41244 31666 41300 31724
rect 41804 31714 41860 31724
rect 41244 31614 41246 31666
rect 41298 31614 41300 31666
rect 41244 28644 41300 31614
rect 41356 31556 41412 31566
rect 41356 31462 41412 31500
rect 41580 30884 41636 30894
rect 41580 30790 41636 30828
rect 41244 28578 41300 28588
rect 41356 30212 41412 30222
rect 41356 28530 41412 30156
rect 41356 28478 41358 28530
rect 41410 28478 41412 28530
rect 41356 28466 41412 28478
rect 41692 28420 41748 28430
rect 41580 26404 41636 26414
rect 41580 26310 41636 26348
rect 41692 20188 41748 28364
rect 41916 26516 41972 31892
rect 42140 31556 42196 32510
rect 42140 31490 42196 31500
rect 42252 28642 42308 28654
rect 42252 28590 42254 28642
rect 42306 28590 42308 28642
rect 42252 28420 42308 28590
rect 42252 28354 42308 28364
rect 41916 26290 41972 26460
rect 42028 26964 42084 26974
rect 42028 26514 42084 26908
rect 42028 26462 42030 26514
rect 42082 26462 42084 26514
rect 42028 26450 42084 26462
rect 41916 26238 41918 26290
rect 41970 26238 41972 26290
rect 41916 26226 41972 26238
rect 42140 26290 42196 26302
rect 42140 26238 42142 26290
rect 42194 26238 42196 26290
rect 42140 26068 42196 26238
rect 42364 26068 42420 26078
rect 42140 26066 42420 26068
rect 42140 26014 42366 26066
rect 42418 26014 42420 26066
rect 42140 26012 42420 26014
rect 42140 20188 42196 26012
rect 42364 26002 42420 26012
rect 41692 20132 41860 20188
rect 42140 20132 42420 20188
rect 41132 17490 41188 17500
rect 41804 3668 41860 20132
rect 41804 3612 42084 3668
rect 41468 3444 41524 3454
rect 41916 3444 41972 3454
rect 41468 3442 41972 3444
rect 41468 3390 41470 3442
rect 41522 3390 41918 3442
rect 41970 3390 41972 3442
rect 41468 3388 41972 3390
rect 41468 3378 41524 3388
rect 40684 3154 40740 3164
rect 41580 800 41636 3388
rect 41916 3378 41972 3388
rect 42028 3332 42084 3612
rect 42252 3332 42308 3342
rect 42028 3330 42308 3332
rect 42028 3278 42254 3330
rect 42306 3278 42308 3330
rect 42028 3276 42308 3278
rect 42252 3266 42308 3276
rect 42364 3332 42420 20132
rect 42476 3556 42532 33404
rect 42700 32676 42756 34972
rect 43148 35028 43204 36540
rect 43484 36594 43540 37436
rect 43484 36542 43486 36594
rect 43538 36542 43540 36594
rect 43484 36530 43540 36542
rect 43708 36484 43764 38668
rect 44604 38724 44660 38734
rect 44604 38630 44660 38668
rect 43708 36418 43764 36428
rect 44716 35922 44772 39004
rect 45276 38994 45332 39004
rect 45500 39060 45556 39340
rect 45500 38928 45556 39004
rect 45612 42532 45668 42590
rect 46060 42532 46116 42542
rect 45612 42530 46116 42532
rect 45612 42478 46062 42530
rect 46114 42478 46116 42530
rect 45612 42476 46116 42478
rect 45612 42084 45668 42476
rect 46060 42466 46116 42476
rect 45388 38836 45444 38846
rect 45388 38742 45444 38780
rect 44716 35870 44718 35922
rect 44770 35870 44772 35922
rect 44716 35812 44772 35870
rect 44716 35746 44772 35756
rect 45164 36484 45220 36494
rect 45164 35922 45220 36428
rect 45164 35870 45166 35922
rect 45218 35870 45220 35922
rect 45164 35700 45220 35870
rect 45164 35634 45220 35644
rect 43148 34962 43204 34972
rect 44716 35028 44772 35038
rect 44716 34934 44772 34972
rect 45164 35028 45220 35038
rect 45164 34356 45220 34972
rect 45164 34224 45220 34300
rect 42700 32544 42756 32620
rect 42700 26516 42756 26526
rect 42700 26422 42756 26460
rect 43036 26178 43092 26190
rect 43036 26126 43038 26178
rect 43090 26126 43092 26178
rect 43036 26066 43092 26126
rect 43036 26014 43038 26066
rect 43090 26014 43092 26066
rect 43036 26002 43092 26014
rect 44268 3668 44324 3678
rect 44268 3574 44324 3612
rect 45164 3666 45220 3678
rect 45164 3614 45166 3666
rect 45218 3614 45220 3666
rect 42476 3490 42532 3500
rect 42364 3266 42420 3276
rect 44492 812 44660 868
rect 44492 800 44548 812
rect 29484 728 29736 800
rect 26824 200 27048 728
rect 29512 200 29736 728
rect 32200 728 32452 800
rect 35560 728 35812 800
rect 32200 200 32424 728
rect 35560 200 35784 728
rect 38248 200 38472 800
rect 41580 728 41832 800
rect 41608 200 41832 728
rect 44296 728 44548 800
rect 44604 756 44660 812
rect 45164 756 45220 3614
rect 45612 3668 45668 42028
rect 48972 40964 49028 40974
rect 47628 40514 47684 40526
rect 47628 40462 47630 40514
rect 47682 40462 47684 40514
rect 47516 40402 47572 40414
rect 47516 40350 47518 40402
rect 47570 40350 47572 40402
rect 47516 39620 47572 40350
rect 47516 39526 47572 39564
rect 47628 40292 47684 40462
rect 47852 40404 47908 40414
rect 47852 40402 48132 40404
rect 47852 40350 47854 40402
rect 47906 40350 48132 40402
rect 47852 40348 48132 40350
rect 47852 40338 47908 40348
rect 46732 39508 46788 39518
rect 46732 39396 46788 39452
rect 47292 39508 47348 39518
rect 47292 39414 47348 39452
rect 47628 39508 47684 40236
rect 48076 39844 48132 40348
rect 48188 40292 48244 40302
rect 48188 40198 48244 40236
rect 48076 39788 48356 39844
rect 48300 39618 48356 39788
rect 48300 39566 48302 39618
rect 48354 39566 48356 39618
rect 48300 39554 48356 39566
rect 47628 39442 47684 39452
rect 47852 39508 47908 39518
rect 46620 39394 46788 39396
rect 46620 39342 46734 39394
rect 46786 39342 46788 39394
rect 46620 39340 46788 39342
rect 46620 39060 46676 39340
rect 46732 39330 46788 39340
rect 47852 39394 47908 39452
rect 48748 39508 48804 39518
rect 48748 39414 48804 39452
rect 48972 39506 49028 40908
rect 48972 39454 48974 39506
rect 49026 39454 49028 39506
rect 47852 39342 47854 39394
rect 47906 39342 47908 39394
rect 47852 39330 47908 39342
rect 48524 39394 48580 39406
rect 48524 39342 48526 39394
rect 48578 39342 48580 39394
rect 46620 38966 46676 39004
rect 45948 38836 46004 38846
rect 45948 38742 46004 38780
rect 48524 38836 48580 39342
rect 48972 39396 49028 39454
rect 49644 39508 49700 39518
rect 49420 39396 49476 39406
rect 48972 39394 49476 39396
rect 48972 39342 49422 39394
rect 49474 39342 49476 39394
rect 48972 39340 49476 39342
rect 48524 38770 48580 38780
rect 45724 38724 45780 38734
rect 45724 38630 45780 38668
rect 46172 38610 46228 38622
rect 46172 38558 46174 38610
rect 46226 38558 46228 38610
rect 46060 36932 46116 36942
rect 45948 35924 46004 35934
rect 45948 35830 46004 35868
rect 46060 35922 46116 36876
rect 46060 35870 46062 35922
rect 46114 35870 46116 35922
rect 45836 35812 45892 35822
rect 45836 35718 45892 35756
rect 46060 35812 46116 35870
rect 46060 35746 46116 35756
rect 46060 35028 46116 35038
rect 46172 35028 46228 38558
rect 49420 36484 49476 39340
rect 49644 37266 49700 39452
rect 49644 37214 49646 37266
rect 49698 37214 49700 37266
rect 49644 37202 49700 37214
rect 49980 37266 50036 37278
rect 49980 37214 49982 37266
rect 50034 37214 50036 37266
rect 49532 37154 49588 37166
rect 49532 37102 49534 37154
rect 49586 37102 49588 37154
rect 49532 36706 49588 37102
rect 49980 37044 50036 37214
rect 49980 36978 50036 36988
rect 49532 36654 49534 36706
rect 49586 36654 49588 36706
rect 49532 36642 49588 36654
rect 49420 36428 49588 36484
rect 49308 36258 49364 36270
rect 49308 36206 49310 36258
rect 49362 36206 49364 36258
rect 47292 35812 47348 35822
rect 47292 35718 47348 35756
rect 46284 35700 46340 35710
rect 46284 35606 46340 35644
rect 46508 35700 46564 35710
rect 46508 35606 46564 35644
rect 46060 35026 46228 35028
rect 46060 34974 46062 35026
rect 46114 34974 46228 35026
rect 46060 34972 46228 34974
rect 46732 35474 46788 35486
rect 46732 35422 46734 35474
rect 46786 35422 46788 35474
rect 46060 34962 46116 34972
rect 45836 34914 45892 34926
rect 45836 34862 45838 34914
rect 45890 34862 45892 34914
rect 45836 34356 45892 34862
rect 46172 34802 46228 34814
rect 46172 34750 46174 34802
rect 46226 34750 46228 34802
rect 46172 34692 46228 34750
rect 46620 34692 46676 34702
rect 46172 34690 46676 34692
rect 46172 34638 46622 34690
rect 46674 34638 46676 34690
rect 46172 34636 46676 34638
rect 45836 34262 45892 34300
rect 45948 34468 46004 34478
rect 45948 34354 46004 34412
rect 45948 34302 45950 34354
rect 46002 34302 46004 34354
rect 45948 34290 46004 34302
rect 46060 33908 46116 33918
rect 46284 33908 46340 33918
rect 46060 33906 46340 33908
rect 46060 33854 46062 33906
rect 46114 33854 46286 33906
rect 46338 33854 46340 33906
rect 46060 33852 46340 33854
rect 46060 33842 46116 33852
rect 46284 33842 46340 33852
rect 46508 20692 46564 34636
rect 46620 34626 46676 34636
rect 46732 34468 46788 35422
rect 49308 35252 49364 36206
rect 49420 36258 49476 36270
rect 49420 36206 49422 36258
rect 49474 36206 49476 36258
rect 49420 35700 49476 36206
rect 49532 35810 49588 36428
rect 49532 35758 49534 35810
rect 49586 35758 49588 35810
rect 49532 35746 49588 35758
rect 49980 36258 50036 36270
rect 49980 36206 49982 36258
rect 50034 36206 50036 36258
rect 49420 35634 49476 35644
rect 49308 35186 49364 35196
rect 49532 35252 49588 35262
rect 46732 34402 46788 34412
rect 46620 34020 46676 34030
rect 46620 34018 46788 34020
rect 46620 33966 46622 34018
rect 46674 33966 46788 34018
rect 46620 33964 46788 33966
rect 46620 33906 46676 33964
rect 46620 33854 46622 33906
rect 46674 33854 46676 33906
rect 46620 33842 46676 33854
rect 46732 23268 46788 33964
rect 49532 33458 49588 35196
rect 49980 35252 50036 36206
rect 49980 35186 50036 35196
rect 50092 35700 50148 46508
rect 52892 46116 52948 46126
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50876 40628 50932 40638
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50764 38948 50820 38958
rect 50876 38948 50932 40572
rect 51324 38948 51380 38958
rect 50764 38946 51380 38948
rect 50764 38894 50766 38946
rect 50818 38894 51326 38946
rect 51378 38894 51380 38946
rect 50764 38892 51380 38894
rect 50764 38882 50820 38892
rect 50876 38610 50932 38622
rect 50876 38558 50878 38610
rect 50930 38558 50932 38610
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50876 37156 50932 38558
rect 50988 37156 51044 37166
rect 50876 37154 51044 37156
rect 50876 37102 50990 37154
rect 51042 37102 51044 37154
rect 50876 37100 51044 37102
rect 50988 37044 51044 37100
rect 50988 36978 51044 36988
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50092 34692 50148 35644
rect 50876 35700 50932 35710
rect 50876 35606 50932 35644
rect 50316 34692 50372 34702
rect 50092 34690 50372 34692
rect 50092 34638 50318 34690
rect 50370 34638 50372 34690
rect 50092 34636 50372 34638
rect 49532 33406 49534 33458
rect 49586 33406 49588 33458
rect 49532 33394 49588 33406
rect 50092 33124 50148 33134
rect 50092 33030 50148 33068
rect 50316 33124 50372 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 33058 50372 33068
rect 50540 33124 50596 33162
rect 50540 33058 50596 33068
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51212 31948 51268 38892
rect 51324 38882 51380 38892
rect 51884 35700 51940 35710
rect 51884 35606 51940 35644
rect 51324 35586 51380 35598
rect 51324 35534 51326 35586
rect 51378 35534 51380 35586
rect 51324 35476 51380 35534
rect 51324 35410 51380 35420
rect 52892 35028 52948 46060
rect 57260 44098 57316 44110
rect 57260 44046 57262 44098
rect 57314 44046 57316 44098
rect 57260 43876 57316 44046
rect 57260 43810 57316 43820
rect 57596 42868 57652 50316
rect 57708 50306 57764 50316
rect 58044 44210 58100 44222
rect 58044 44158 58046 44210
rect 58098 44158 58100 44210
rect 57596 42802 57652 42812
rect 57708 44098 57764 44110
rect 57708 44046 57710 44098
rect 57762 44046 57764 44098
rect 57708 41188 57764 44046
rect 58044 43876 58100 44158
rect 58044 43810 58100 43820
rect 57596 41132 57764 41188
rect 57260 41076 57316 41086
rect 57260 40982 57316 41020
rect 57596 37940 57652 41132
rect 58044 41076 58100 41086
rect 58044 40982 58100 41020
rect 57708 40962 57764 40974
rect 57708 40910 57710 40962
rect 57762 40910 57764 40962
rect 57708 40404 57764 40910
rect 57708 40338 57764 40348
rect 57596 37874 57652 37884
rect 58044 37938 58100 37950
rect 58044 37886 58046 37938
rect 58098 37886 58100 37938
rect 57260 37828 57316 37838
rect 57260 37734 57316 37772
rect 57708 37826 57764 37838
rect 57708 37774 57710 37826
rect 57762 37774 57764 37826
rect 57708 37492 57764 37774
rect 58044 37828 58100 37886
rect 58044 37762 58100 37772
rect 57708 37426 57764 37436
rect 52892 34962 52948 34972
rect 56252 35028 56308 35038
rect 56252 34934 56308 34972
rect 56812 35028 56868 35038
rect 56812 34914 56868 34972
rect 57820 35028 57876 35038
rect 57820 34934 57876 34972
rect 56812 34862 56814 34914
rect 56866 34862 56868 34914
rect 56812 34850 56868 34862
rect 57708 33124 57764 33134
rect 51212 31892 51380 31948
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 46732 23202 46788 23212
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 46508 20626 46564 20636
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 51324 14644 51380 31892
rect 57484 31220 57540 31230
rect 56252 27748 56308 27758
rect 56252 25620 56308 27692
rect 56252 25618 56868 25620
rect 56252 25566 56254 25618
rect 56306 25566 56868 25618
rect 56252 25564 56868 25566
rect 56252 25554 56308 25564
rect 56812 25506 56868 25564
rect 56812 25454 56814 25506
rect 56866 25454 56868 25506
rect 56812 25442 56868 25454
rect 57260 20578 57316 20590
rect 57260 20526 57262 20578
rect 57314 20526 57316 20578
rect 57260 20356 57316 20526
rect 57260 20290 57316 20300
rect 57260 17444 57316 17454
rect 57260 17350 57316 17388
rect 51324 14578 51380 14588
rect 56364 14644 56420 14654
rect 56364 14550 56420 14588
rect 56812 14644 56868 14654
rect 56812 14530 56868 14588
rect 56812 14478 56814 14530
rect 56866 14478 56868 14530
rect 56812 14466 56868 14478
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 56812 11394 56868 11406
rect 56812 11342 56814 11394
rect 56866 11342 56868 11394
rect 56364 11172 56420 11182
rect 56364 11078 56420 11116
rect 56812 11172 56868 11342
rect 56812 11106 56868 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 57484 8428 57540 31164
rect 57596 30884 57652 30894
rect 57596 20188 57652 30828
rect 57708 29650 57764 33068
rect 58044 31556 58100 31566
rect 58044 31462 58100 31500
rect 57708 29598 57710 29650
rect 57762 29598 57764 29650
rect 57708 29586 57764 29598
rect 58044 29428 58100 29438
rect 58044 29426 58212 29428
rect 58044 29374 58046 29426
rect 58098 29374 58212 29426
rect 58044 29372 58212 29374
rect 58044 29362 58100 29372
rect 58156 28868 58212 29372
rect 58156 28754 58212 28812
rect 58156 28702 58158 28754
rect 58210 28702 58212 28754
rect 58156 28690 58212 28702
rect 57820 25620 57876 25630
rect 57820 25526 57876 25564
rect 57708 23268 57764 23278
rect 57708 23174 57764 23212
rect 58044 23154 58100 23166
rect 58044 23102 58046 23154
rect 58098 23102 58100 23154
rect 58044 23044 58100 23102
rect 58044 22484 58100 22988
rect 58156 22484 58212 22494
rect 58044 22482 58212 22484
rect 58044 22430 58158 22482
rect 58210 22430 58212 22482
rect 58044 22428 58212 22430
rect 58156 22418 58212 22428
rect 57708 20692 57764 20702
rect 57708 20598 57764 20636
rect 58044 20690 58100 20702
rect 58044 20638 58046 20690
rect 58098 20638 58100 20690
rect 58044 20356 58100 20638
rect 58044 20290 58100 20300
rect 57596 20132 57876 20188
rect 57708 17556 57764 17566
rect 57708 17462 57764 17500
rect 57708 14418 57764 14430
rect 57708 14366 57710 14418
rect 57762 14366 57764 14418
rect 57708 14308 57764 14366
rect 57708 14242 57764 14252
rect 57708 11282 57764 11294
rect 57708 11230 57710 11282
rect 57762 11230 57764 11282
rect 57708 10948 57764 11230
rect 57708 10882 57764 10892
rect 57484 8372 57652 8428
rect 57260 8036 57316 8046
rect 57260 7942 57316 7980
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 57260 5012 57316 5022
rect 57596 5012 57652 8372
rect 57708 8148 57764 8158
rect 57708 8054 57764 8092
rect 57708 5012 57764 5022
rect 57596 5010 57764 5012
rect 57596 4958 57710 5010
rect 57762 4958 57764 5010
rect 57596 4956 57764 4958
rect 57260 4918 57316 4956
rect 57708 4946 57764 4956
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 57708 4564 57764 4574
rect 57820 4564 57876 20132
rect 58044 17554 58100 17566
rect 58044 17502 58046 17554
rect 58098 17502 58100 17554
rect 58044 17444 58100 17502
rect 58044 16996 58100 17388
rect 58044 16930 58100 16940
rect 58044 8148 58100 8158
rect 58044 8054 58100 8092
rect 58044 6018 58100 6030
rect 58044 5966 58046 6018
rect 58098 5966 58100 6018
rect 58044 5236 58100 5966
rect 58044 5170 58100 5180
rect 58044 5012 58100 5022
rect 58100 4956 58212 5012
rect 58044 4880 58100 4956
rect 57708 4562 57876 4564
rect 57708 4510 57710 4562
rect 57762 4510 57876 4562
rect 57708 4508 57876 4510
rect 57708 4498 57764 4508
rect 58044 4338 58100 4350
rect 58044 4286 58046 4338
rect 58098 4286 58100 4338
rect 56812 4228 56868 4238
rect 56812 4134 56868 4172
rect 58044 4228 58100 4286
rect 45612 3556 45668 3612
rect 45948 3556 46004 3566
rect 45612 3554 46004 3556
rect 45612 3502 45950 3554
rect 46002 3502 46004 3554
rect 45612 3500 46004 3502
rect 45948 3490 46004 3500
rect 56028 3556 56084 3566
rect 56028 3462 56084 3500
rect 56700 3556 56756 3566
rect 56700 3462 56756 3500
rect 48188 3444 48244 3454
rect 47852 812 48020 868
rect 47852 800 47908 812
rect 44296 200 44520 728
rect 44604 700 45220 756
rect 47656 728 47908 800
rect 47964 756 48020 812
rect 48188 756 48244 3388
rect 49196 3444 49252 3454
rect 49196 3350 49252 3388
rect 50204 3444 50260 3454
rect 50428 3444 50484 3454
rect 50204 3442 50428 3444
rect 50204 3390 50206 3442
rect 50258 3390 50428 3442
rect 50204 3388 50428 3390
rect 50204 3378 50260 3388
rect 48860 3330 48916 3342
rect 48860 3278 48862 3330
rect 48914 3278 48916 3330
rect 48860 3220 48916 3278
rect 48860 3154 48916 3164
rect 50428 800 50484 3388
rect 50988 3444 51044 3454
rect 50652 3332 50708 3370
rect 50988 3350 51044 3388
rect 56588 3444 56644 3454
rect 50652 3266 50708 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 56588 800 56644 3388
rect 57596 3444 57652 3454
rect 57596 3350 57652 3388
rect 58044 2884 58100 4172
rect 58044 2818 58100 2828
rect 47656 200 47880 728
rect 47964 700 48244 756
rect 50344 200 50568 800
rect 53704 200 53928 800
rect 56392 728 56644 800
rect 58156 756 58212 4956
rect 58940 812 59108 868
rect 58940 756 58996 812
rect 56392 200 56616 728
rect 58156 700 58996 756
rect 59052 800 59108 812
rect 59052 728 59304 800
rect 59080 200 59304 728
<< via2 >>
rect 1820 56364 1876 56420
rect 4844 56140 4900 56196
rect 6076 56194 6132 56196
rect 6076 56142 6078 56194
rect 6078 56142 6130 56194
rect 6130 56142 6132 56194
rect 6076 56140 6132 56142
rect 3500 55916 3556 55972
rect 4060 55970 4116 55972
rect 4060 55918 4062 55970
rect 4062 55918 4114 55970
rect 4114 55918 4116 55970
rect 4060 55916 4116 55918
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 2044 53788 2100 53844
rect 1820 53170 1876 53172
rect 1820 53118 1822 53170
rect 1822 53118 1874 53170
rect 1874 53118 1876 53170
rect 1820 53116 1876 53118
rect 1820 50482 1876 50484
rect 1820 50430 1822 50482
rect 1822 50430 1874 50482
rect 1874 50430 1876 50482
rect 1820 50428 1876 50430
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 3724 53842 3780 53844
rect 3724 53790 3726 53842
rect 3726 53790 3778 53842
rect 3778 53790 3780 53842
rect 3724 53788 3780 53790
rect 2268 53004 2324 53060
rect 2156 51436 2212 51492
rect 3388 51100 3444 51156
rect 2156 48748 2212 48804
rect 2044 47852 2100 47908
rect 2044 47068 2100 47124
rect 1820 44434 1876 44436
rect 1820 44382 1822 44434
rect 1822 44382 1874 44434
rect 1874 44382 1876 44434
rect 1820 44380 1876 44382
rect 2492 46508 2548 46564
rect 3164 46562 3220 46564
rect 3164 46510 3166 46562
rect 3166 46510 3218 46562
rect 3218 46510 3220 46562
rect 3164 46508 3220 46510
rect 3276 45612 3332 45668
rect 1820 41804 1876 41860
rect 1820 38220 1876 38276
rect 1708 35810 1764 35812
rect 1708 35758 1710 35810
rect 1710 35758 1762 35810
rect 1762 35758 1764 35810
rect 1708 35756 1764 35758
rect 3724 53058 3780 53060
rect 3724 53006 3726 53058
rect 3726 53006 3778 53058
rect 3778 53006 3780 53058
rect 3724 53004 3780 53006
rect 3724 48748 3780 48804
rect 3948 52780 4004 52836
rect 3948 50316 4004 50372
rect 4060 48972 4116 49028
rect 6188 53058 6244 53060
rect 6188 53006 6190 53058
rect 6190 53006 6242 53058
rect 6242 53006 6244 53058
rect 6188 53004 6244 53006
rect 4508 52834 4564 52836
rect 4508 52782 4510 52834
rect 4510 52782 4562 52834
rect 4562 52782 4564 52834
rect 4508 52780 4564 52782
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4620 51490 4676 51492
rect 4620 51438 4622 51490
rect 4622 51438 4674 51490
rect 4674 51438 4676 51490
rect 4620 51436 4676 51438
rect 4732 51154 4788 51156
rect 4732 51102 4734 51154
rect 4734 51102 4786 51154
rect 4786 51102 4788 51154
rect 4732 51100 4788 51102
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 5180 50316 5236 50372
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4956 48972 5012 49028
rect 4508 48748 4564 48804
rect 3948 48354 4004 48356
rect 3948 48302 3950 48354
rect 3950 48302 4002 48354
rect 4002 48302 4004 48354
rect 3948 48300 4004 48302
rect 3836 47292 3892 47348
rect 3724 47068 3780 47124
rect 3724 46674 3780 46676
rect 3724 46622 3726 46674
rect 3726 46622 3778 46674
rect 3778 46622 3780 46674
rect 3724 46620 3780 46622
rect 4508 48300 4564 48356
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4844 47292 4900 47348
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 3948 39452 4004 39508
rect 4172 42588 4228 42644
rect 3612 36652 3668 36708
rect 3836 38722 3892 38724
rect 3836 38670 3838 38722
rect 3838 38670 3890 38722
rect 3890 38670 3892 38722
rect 3836 38668 3892 38670
rect 3500 36428 3556 36484
rect 3388 35868 3444 35924
rect 2156 34188 2212 34244
rect 3500 35420 3556 35476
rect 2044 32450 2100 32452
rect 2044 32398 2046 32450
rect 2046 32398 2098 32450
rect 2098 32398 2100 32450
rect 2044 32396 2100 32398
rect 2268 30828 2324 30884
rect 2156 30268 2212 30324
rect 1820 29650 1876 29652
rect 1820 29598 1822 29650
rect 1822 29598 1874 29650
rect 1874 29598 1876 29650
rect 1820 29596 1876 29598
rect 2156 26348 2212 26404
rect 2156 23660 2212 23716
rect 2044 20972 2100 21028
rect 2156 18620 2212 18676
rect 1820 17554 1876 17556
rect 1820 17502 1822 17554
rect 1822 17502 1874 17554
rect 1874 17502 1876 17554
rect 1820 17500 1876 17502
rect 3948 38610 4004 38612
rect 3948 38558 3950 38610
rect 3950 38558 4002 38610
rect 4002 38558 4004 38610
rect 3948 38556 4004 38558
rect 3836 36706 3892 36708
rect 3836 36654 3838 36706
rect 3838 36654 3890 36706
rect 3890 36654 3892 36706
rect 3836 36652 3892 36654
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5180 48748 5236 48804
rect 5404 47516 5460 47572
rect 5852 47516 5908 47572
rect 4844 39004 4900 39060
rect 4396 38722 4452 38724
rect 4396 38670 4398 38722
rect 4398 38670 4450 38722
rect 4450 38670 4452 38722
rect 4396 38668 4452 38670
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 5068 38444 5124 38500
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4060 36594 4116 36596
rect 4060 36542 4062 36594
rect 4062 36542 4114 36594
rect 4114 36542 4116 36594
rect 4060 36540 4116 36542
rect 4396 36316 4452 36372
rect 4508 36258 4564 36260
rect 4508 36206 4510 36258
rect 4510 36206 4562 36258
rect 4562 36206 4564 36258
rect 4508 36204 4564 36206
rect 4732 35980 4788 36036
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5068 36316 5124 36372
rect 5292 35980 5348 36036
rect 4732 34242 4788 34244
rect 4732 34190 4734 34242
rect 4734 34190 4786 34242
rect 4786 34190 4788 34242
rect 4732 34188 4788 34190
rect 5628 36652 5684 36708
rect 5516 35308 5572 35364
rect 4956 34018 5012 34020
rect 4956 33966 4958 34018
rect 4958 33966 5010 34018
rect 5010 33966 5012 34018
rect 4956 33964 5012 33966
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5628 31836 5684 31892
rect 5516 30994 5572 30996
rect 5516 30942 5518 30994
rect 5518 30942 5570 30994
rect 5570 30942 5572 30994
rect 5516 30940 5572 30942
rect 4732 30882 4788 30884
rect 4732 30830 4734 30882
rect 4734 30830 4786 30882
rect 4786 30830 4788 30882
rect 4732 30828 4788 30830
rect 5180 30882 5236 30884
rect 5180 30830 5182 30882
rect 5182 30830 5234 30882
rect 5234 30830 5236 30882
rect 5180 30828 5236 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5516 30380 5572 30436
rect 5740 30322 5796 30324
rect 5740 30270 5742 30322
rect 5742 30270 5794 30322
rect 5794 30270 5796 30322
rect 5740 30268 5796 30270
rect 6188 45218 6244 45220
rect 6188 45166 6190 45218
rect 6190 45166 6242 45218
rect 6242 45166 6244 45218
rect 6188 45164 6244 45166
rect 6188 43762 6244 43764
rect 6188 43710 6190 43762
rect 6190 43710 6242 43762
rect 6242 43710 6244 43762
rect 6188 43708 6244 43710
rect 6188 40908 6244 40964
rect 5964 30882 6020 30884
rect 5964 30830 5966 30882
rect 5966 30830 6018 30882
rect 6018 30830 6020 30882
rect 5964 30828 6020 30830
rect 5964 30492 6020 30548
rect 6076 30322 6132 30324
rect 6076 30270 6078 30322
rect 6078 30270 6130 30322
rect 6130 30270 6132 30322
rect 6076 30268 6132 30270
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3052 26908 3108 26964
rect 3500 26908 3556 26964
rect 6076 28082 6132 28084
rect 6076 28030 6078 28082
rect 6078 28030 6130 28082
rect 6130 28030 6132 28082
rect 6076 28028 6132 28030
rect 6076 27746 6132 27748
rect 6076 27694 6078 27746
rect 6078 27694 6130 27746
rect 6130 27694 6132 27746
rect 6076 27692 6132 27694
rect 2380 26572 2436 26628
rect 1820 14700 1876 14756
rect 2044 11564 2100 11620
rect 4284 26012 4340 26068
rect 3052 23996 3108 24052
rect 3612 24050 3668 24052
rect 3612 23998 3614 24050
rect 3614 23998 3666 24050
rect 3666 23998 3668 24050
rect 3612 23996 3668 23998
rect 3500 23660 3556 23716
rect 3612 22316 3668 22372
rect 3052 12348 3108 12404
rect 3500 12402 3556 12404
rect 3500 12350 3502 12402
rect 3502 12350 3554 12402
rect 3554 12350 3556 12402
rect 3500 12348 3556 12350
rect 1820 8652 1876 8708
rect 3948 21756 4004 21812
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5852 23996 5908 24052
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3724 18620 3780 18676
rect 3052 6076 3108 6132
rect 2044 5516 2100 5572
rect 3052 5180 3108 5236
rect 812 4956 868 5012
rect 2156 5010 2212 5012
rect 2156 4958 2158 5010
rect 2158 4958 2210 5010
rect 2210 4958 2212 5010
rect 2156 4956 2212 4958
rect 3500 6130 3556 6132
rect 3500 6078 3502 6130
rect 3502 6078 3554 6130
rect 3554 6078 3556 6130
rect 3500 6076 3556 6078
rect 3612 5234 3668 5236
rect 3612 5182 3614 5234
rect 3614 5182 3666 5234
rect 3666 5182 3668 5234
rect 3612 5180 3668 5182
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 6524 48524 6580 48580
rect 6412 36482 6468 36484
rect 6412 36430 6414 36482
rect 6414 36430 6466 36482
rect 6466 36430 6468 36482
rect 6412 36428 6468 36430
rect 6300 35420 6356 35476
rect 6412 31836 6468 31892
rect 6412 31388 6468 31444
rect 6300 30828 6356 30884
rect 6300 28028 6356 28084
rect 6188 5180 6244 5236
rect 6300 27858 6356 27860
rect 6300 27806 6302 27858
rect 6302 27806 6354 27858
rect 6354 27806 6356 27858
rect 6300 27804 6356 27806
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 2044 2828 2100 2884
rect 6636 42754 6692 42756
rect 6636 42702 6638 42754
rect 6638 42702 6690 42754
rect 6690 42702 6692 42754
rect 6636 42700 6692 42702
rect 6636 40962 6692 40964
rect 6636 40910 6638 40962
rect 6638 40910 6690 40962
rect 6690 40910 6692 40962
rect 6636 40908 6692 40910
rect 6860 35756 6916 35812
rect 6524 30492 6580 30548
rect 6748 27858 6804 27860
rect 6748 27806 6750 27858
rect 6750 27806 6802 27858
rect 6802 27806 6804 27858
rect 6748 27804 6804 27806
rect 7084 42252 7140 42308
rect 7644 55916 7700 55972
rect 8316 55074 8372 55076
rect 8316 55022 8318 55074
rect 8318 55022 8370 55074
rect 8370 55022 8372 55074
rect 8316 55020 8372 55022
rect 10780 55020 10836 55076
rect 11452 54796 11508 54852
rect 11452 54236 11508 54292
rect 8204 52892 8260 52948
rect 7980 51938 8036 51940
rect 7980 51886 7982 51938
rect 7982 51886 8034 51938
rect 8034 51886 8036 51938
rect 7980 51884 8036 51886
rect 7420 48802 7476 48804
rect 7420 48750 7422 48802
rect 7422 48750 7474 48802
rect 7474 48750 7476 48802
rect 7420 48748 7476 48750
rect 7756 45276 7812 45332
rect 7420 40962 7476 40964
rect 7420 40910 7422 40962
rect 7422 40910 7474 40962
rect 7474 40910 7476 40962
rect 7420 40908 7476 40910
rect 7196 39900 7252 39956
rect 7308 36482 7364 36484
rect 7308 36430 7310 36482
rect 7310 36430 7362 36482
rect 7362 36430 7364 36482
rect 7308 36428 7364 36430
rect 7532 36316 7588 36372
rect 7308 28082 7364 28084
rect 7308 28030 7310 28082
rect 7310 28030 7362 28082
rect 7362 28030 7364 28082
rect 7308 28028 7364 28030
rect 9100 53730 9156 53732
rect 9100 53678 9102 53730
rect 9102 53678 9154 53730
rect 9154 53678 9156 53730
rect 9100 53676 9156 53678
rect 12348 55074 12404 55076
rect 12348 55022 12350 55074
rect 12350 55022 12402 55074
rect 12402 55022 12404 55074
rect 12348 55020 12404 55022
rect 12124 53618 12180 53620
rect 12124 53566 12126 53618
rect 12126 53566 12178 53618
rect 12178 53566 12180 53618
rect 12124 53564 12180 53566
rect 11900 53452 11956 53508
rect 11564 53116 11620 53172
rect 12348 53116 12404 53172
rect 12460 53676 12516 53732
rect 10556 53004 10612 53060
rect 8652 52892 8708 52948
rect 9100 52946 9156 52948
rect 9100 52894 9102 52946
rect 9102 52894 9154 52946
rect 9154 52894 9156 52946
rect 9100 52892 9156 52894
rect 9660 52892 9716 52948
rect 8540 52780 8596 52836
rect 10220 52834 10276 52836
rect 10220 52782 10222 52834
rect 10222 52782 10274 52834
rect 10274 52782 10276 52834
rect 10220 52780 10276 52782
rect 9660 52108 9716 52164
rect 10220 52220 10276 52276
rect 10556 52556 10612 52612
rect 11900 52274 11956 52276
rect 11900 52222 11902 52274
rect 11902 52222 11954 52274
rect 11954 52222 11956 52274
rect 11900 52220 11956 52222
rect 10892 52162 10948 52164
rect 10892 52110 10894 52162
rect 10894 52110 10946 52162
rect 10946 52110 10948 52162
rect 10892 52108 10948 52110
rect 11452 52162 11508 52164
rect 11452 52110 11454 52162
rect 11454 52110 11506 52162
rect 11506 52110 11508 52162
rect 11452 52108 11508 52110
rect 11116 51884 11172 51940
rect 11116 51378 11172 51380
rect 11116 51326 11118 51378
rect 11118 51326 11170 51378
rect 11170 51326 11172 51378
rect 11116 51324 11172 51326
rect 10332 50764 10388 50820
rect 8652 50428 8708 50484
rect 11228 50428 11284 50484
rect 11004 49868 11060 49924
rect 11116 49532 11172 49588
rect 9772 48748 9828 48804
rect 10556 48860 10612 48916
rect 11452 49868 11508 49924
rect 11340 48802 11396 48804
rect 11340 48750 11342 48802
rect 11342 48750 11394 48802
rect 11394 48750 11396 48802
rect 11340 48748 11396 48750
rect 8540 45106 8596 45108
rect 8540 45054 8542 45106
rect 8542 45054 8594 45106
rect 8594 45054 8596 45106
rect 8540 45052 8596 45054
rect 9100 46508 9156 46564
rect 7980 36764 8036 36820
rect 8092 44044 8148 44100
rect 8204 43260 8260 43316
rect 8540 43148 8596 43204
rect 10668 45948 10724 46004
rect 10108 45890 10164 45892
rect 10108 45838 10110 45890
rect 10110 45838 10162 45890
rect 10162 45838 10164 45890
rect 10108 45836 10164 45838
rect 11228 46002 11284 46004
rect 11228 45950 11230 46002
rect 11230 45950 11282 46002
rect 11282 45950 11284 46002
rect 11228 45948 11284 45950
rect 9884 45164 9940 45220
rect 9436 45052 9492 45108
rect 8876 43372 8932 43428
rect 8876 42700 8932 42756
rect 8204 38556 8260 38612
rect 8988 36652 9044 36708
rect 8876 36594 8932 36596
rect 8876 36542 8878 36594
rect 8878 36542 8930 36594
rect 8930 36542 8932 36594
rect 8876 36540 8932 36542
rect 8652 36316 8708 36372
rect 8204 35922 8260 35924
rect 8204 35870 8206 35922
rect 8206 35870 8258 35922
rect 8258 35870 8260 35922
rect 8204 35868 8260 35870
rect 7980 35756 8036 35812
rect 8540 35084 8596 35140
rect 7980 34300 8036 34356
rect 8540 34354 8596 34356
rect 8540 34302 8542 34354
rect 8542 34302 8594 34354
rect 8594 34302 8596 34354
rect 8540 34300 8596 34302
rect 8092 34242 8148 34244
rect 8092 34190 8094 34242
rect 8094 34190 8146 34242
rect 8146 34190 8148 34242
rect 8092 34188 8148 34190
rect 8764 36204 8820 36260
rect 9212 36204 9268 36260
rect 9212 35756 9268 35812
rect 8988 35308 9044 35364
rect 9100 34748 9156 34804
rect 8876 34188 8932 34244
rect 8652 33852 8708 33908
rect 7868 32060 7924 32116
rect 8652 33292 8708 33348
rect 8540 31276 8596 31332
rect 8540 30492 8596 30548
rect 7644 27244 7700 27300
rect 9772 44716 9828 44772
rect 9772 43708 9828 43764
rect 9548 43596 9604 43652
rect 9660 43426 9716 43428
rect 9660 43374 9662 43426
rect 9662 43374 9714 43426
rect 9714 43374 9716 43426
rect 9660 43372 9716 43374
rect 10780 45276 10836 45332
rect 10780 44828 10836 44884
rect 10556 44322 10612 44324
rect 10556 44270 10558 44322
rect 10558 44270 10610 44322
rect 10610 44270 10612 44322
rect 10556 44268 10612 44270
rect 11228 45106 11284 45108
rect 11228 45054 11230 45106
rect 11230 45054 11282 45106
rect 11282 45054 11284 45106
rect 11228 45052 11284 45054
rect 10220 43650 10276 43652
rect 10220 43598 10222 43650
rect 10222 43598 10274 43650
rect 10274 43598 10276 43650
rect 10220 43596 10276 43598
rect 10108 43372 10164 43428
rect 10668 43372 10724 43428
rect 9884 43036 9940 43092
rect 11452 48412 11508 48468
rect 11116 43372 11172 43428
rect 10780 43148 10836 43204
rect 9772 41020 9828 41076
rect 10108 36258 10164 36260
rect 10108 36206 10110 36258
rect 10110 36206 10162 36258
rect 10162 36206 10164 36258
rect 10108 36204 10164 36206
rect 9772 35810 9828 35812
rect 9772 35758 9774 35810
rect 9774 35758 9826 35810
rect 9826 35758 9828 35810
rect 9772 35756 9828 35758
rect 9884 35980 9940 36036
rect 9436 33740 9492 33796
rect 9548 35308 9604 35364
rect 9212 30434 9268 30436
rect 9212 30382 9214 30434
rect 9214 30382 9266 30434
rect 9266 30382 9268 30434
rect 9212 30380 9268 30382
rect 6860 23660 6916 23716
rect 9436 30604 9492 30660
rect 9436 30434 9492 30436
rect 9436 30382 9438 30434
rect 9438 30382 9490 30434
rect 9490 30382 9492 30434
rect 9436 30380 9492 30382
rect 9324 29260 9380 29316
rect 10108 35868 10164 35924
rect 11116 42252 11172 42308
rect 10556 40908 10612 40964
rect 10556 40514 10612 40516
rect 10556 40462 10558 40514
rect 10558 40462 10610 40514
rect 10610 40462 10612 40514
rect 10556 40460 10612 40462
rect 10892 38444 10948 38500
rect 10892 37212 10948 37268
rect 10444 35420 10500 35476
rect 9884 34076 9940 34132
rect 9772 34018 9828 34020
rect 9772 33966 9774 34018
rect 9774 33966 9826 34018
rect 9826 33966 9828 34018
rect 9772 33964 9828 33966
rect 9660 32956 9716 33012
rect 9996 34636 10052 34692
rect 9996 33740 10052 33796
rect 10220 34802 10276 34804
rect 10220 34750 10222 34802
rect 10222 34750 10274 34802
rect 10274 34750 10276 34802
rect 10220 34748 10276 34750
rect 10332 34690 10388 34692
rect 10332 34638 10334 34690
rect 10334 34638 10386 34690
rect 10386 34638 10388 34690
rect 10332 34636 10388 34638
rect 10556 34354 10612 34356
rect 10556 34302 10558 34354
rect 10558 34302 10610 34354
rect 10610 34302 10612 34354
rect 10556 34300 10612 34302
rect 10780 34802 10836 34804
rect 10780 34750 10782 34802
rect 10782 34750 10834 34802
rect 10834 34750 10836 34802
rect 10780 34748 10836 34750
rect 10444 34242 10500 34244
rect 10444 34190 10446 34242
rect 10446 34190 10498 34242
rect 10498 34190 10500 34242
rect 10444 34188 10500 34190
rect 10668 34130 10724 34132
rect 10668 34078 10670 34130
rect 10670 34078 10722 34130
rect 10722 34078 10724 34130
rect 10668 34076 10724 34078
rect 10220 33852 10276 33908
rect 10108 32562 10164 32564
rect 10108 32510 10110 32562
rect 10110 32510 10162 32562
rect 10162 32510 10164 32562
rect 10108 32508 10164 32510
rect 9772 32060 9828 32116
rect 9660 30492 9716 30548
rect 9660 29484 9716 29540
rect 7756 26572 7812 26628
rect 9996 30604 10052 30660
rect 9884 30210 9940 30212
rect 9884 30158 9886 30210
rect 9886 30158 9938 30210
rect 9938 30158 9940 30210
rect 9884 30156 9940 30158
rect 10108 30098 10164 30100
rect 10108 30046 10110 30098
rect 10110 30046 10162 30098
rect 10162 30046 10164 30098
rect 10108 30044 10164 30046
rect 10108 27746 10164 27748
rect 10108 27694 10110 27746
rect 10110 27694 10162 27746
rect 10162 27694 10164 27746
rect 10108 27692 10164 27694
rect 10444 31836 10500 31892
rect 10444 30492 10500 30548
rect 10332 30044 10388 30100
rect 10780 33516 10836 33572
rect 10892 32620 10948 32676
rect 11004 32060 11060 32116
rect 11004 31890 11060 31892
rect 11004 31838 11006 31890
rect 11006 31838 11058 31890
rect 11058 31838 11060 31890
rect 11004 31836 11060 31838
rect 10892 31218 10948 31220
rect 10892 31166 10894 31218
rect 10894 31166 10946 31218
rect 10946 31166 10948 31218
rect 10892 31164 10948 31166
rect 10668 30044 10724 30100
rect 11004 29596 11060 29652
rect 11340 43260 11396 43316
rect 11340 42924 11396 42980
rect 11340 40962 11396 40964
rect 11340 40910 11342 40962
rect 11342 40910 11394 40962
rect 11394 40910 11396 40962
rect 11340 40908 11396 40910
rect 11340 38332 11396 38388
rect 11452 37154 11508 37156
rect 11452 37102 11454 37154
rect 11454 37102 11506 37154
rect 11506 37102 11508 37154
rect 11452 37100 11508 37102
rect 11452 36428 11508 36484
rect 11340 35420 11396 35476
rect 11228 34300 11284 34356
rect 11340 35084 11396 35140
rect 11228 34130 11284 34132
rect 11228 34078 11230 34130
rect 11230 34078 11282 34130
rect 11282 34078 11284 34130
rect 11228 34076 11284 34078
rect 11228 33404 11284 33460
rect 10332 27804 10388 27860
rect 10556 29426 10612 29428
rect 10556 29374 10558 29426
rect 10558 29374 10610 29426
rect 10610 29374 10612 29426
rect 10556 29372 10612 29374
rect 10332 27634 10388 27636
rect 10332 27582 10334 27634
rect 10334 27582 10386 27634
rect 10386 27582 10388 27634
rect 10332 27580 10388 27582
rect 10556 28588 10612 28644
rect 10220 26684 10276 26740
rect 10220 26514 10276 26516
rect 10220 26462 10222 26514
rect 10222 26462 10274 26514
rect 10274 26462 10276 26514
rect 10220 26460 10276 26462
rect 10220 26012 10276 26068
rect 9772 25394 9828 25396
rect 9772 25342 9774 25394
rect 9774 25342 9826 25394
rect 9826 25342 9828 25394
rect 9772 25340 9828 25342
rect 10556 26908 10612 26964
rect 10332 25340 10388 25396
rect 12236 49922 12292 49924
rect 12236 49870 12238 49922
rect 12238 49870 12290 49922
rect 12290 49870 12292 49922
rect 12236 49868 12292 49870
rect 11900 49532 11956 49588
rect 12124 48466 12180 48468
rect 12124 48414 12126 48466
rect 12126 48414 12178 48466
rect 12178 48414 12180 48466
rect 12124 48412 12180 48414
rect 11676 45890 11732 45892
rect 11676 45838 11678 45890
rect 11678 45838 11730 45890
rect 11730 45838 11732 45890
rect 11676 45836 11732 45838
rect 12348 46562 12404 46564
rect 12348 46510 12350 46562
rect 12350 46510 12402 46562
rect 12402 46510 12404 46562
rect 12348 46508 12404 46510
rect 12124 44322 12180 44324
rect 12124 44270 12126 44322
rect 12126 44270 12178 44322
rect 12178 44270 12180 44322
rect 12124 44268 12180 44270
rect 11676 43372 11732 43428
rect 12124 43426 12180 43428
rect 12124 43374 12126 43426
rect 12126 43374 12178 43426
rect 12178 43374 12180 43426
rect 12124 43372 12180 43374
rect 11788 37324 11844 37380
rect 12012 38220 12068 38276
rect 11900 36652 11956 36708
rect 12012 36876 12068 36932
rect 11900 36482 11956 36484
rect 11900 36430 11902 36482
rect 11902 36430 11954 36482
rect 11954 36430 11956 36482
rect 11900 36428 11956 36430
rect 11900 36204 11956 36260
rect 11564 35084 11620 35140
rect 11676 35420 11732 35476
rect 11452 33516 11508 33572
rect 11788 34748 11844 34804
rect 12012 35868 12068 35924
rect 11676 33852 11732 33908
rect 11452 32786 11508 32788
rect 11452 32734 11454 32786
rect 11454 32734 11506 32786
rect 11506 32734 11508 32786
rect 11452 32732 11508 32734
rect 11564 32674 11620 32676
rect 11564 32622 11566 32674
rect 11566 32622 11618 32674
rect 11618 32622 11620 32674
rect 11564 32620 11620 32622
rect 11340 31164 11396 31220
rect 11900 33458 11956 33460
rect 11900 33406 11902 33458
rect 11902 33406 11954 33458
rect 11954 33406 11956 33458
rect 11900 33404 11956 33406
rect 11900 33180 11956 33236
rect 12236 35980 12292 36036
rect 12236 35644 12292 35700
rect 11900 31836 11956 31892
rect 11788 31724 11844 31780
rect 11340 30994 11396 30996
rect 11340 30942 11342 30994
rect 11342 30942 11394 30994
rect 11394 30942 11396 30994
rect 11340 30940 11396 30942
rect 11340 29986 11396 29988
rect 11340 29934 11342 29986
rect 11342 29934 11394 29986
rect 11394 29934 11396 29986
rect 11340 29932 11396 29934
rect 11340 29372 11396 29428
rect 11116 29148 11172 29204
rect 11004 27858 11060 27860
rect 11004 27806 11006 27858
rect 11006 27806 11058 27858
rect 11058 27806 11060 27858
rect 11004 27804 11060 27806
rect 10892 26012 10948 26068
rect 10444 23436 10500 23492
rect 10556 24780 10612 24836
rect 10332 22370 10388 22372
rect 10332 22318 10334 22370
rect 10334 22318 10386 22370
rect 10386 22318 10388 22370
rect 10332 22316 10388 22318
rect 11900 31666 11956 31668
rect 11900 31614 11902 31666
rect 11902 31614 11954 31666
rect 11954 31614 11956 31666
rect 11900 31612 11956 31614
rect 11676 31554 11732 31556
rect 11676 31502 11678 31554
rect 11678 31502 11730 31554
rect 11730 31502 11732 31554
rect 11676 31500 11732 31502
rect 12236 32508 12292 32564
rect 11788 30380 11844 30436
rect 12124 31836 12180 31892
rect 11564 27858 11620 27860
rect 11564 27806 11566 27858
rect 11566 27806 11618 27858
rect 11618 27806 11620 27858
rect 11564 27804 11620 27806
rect 11452 27580 11508 27636
rect 12012 31106 12068 31108
rect 12012 31054 12014 31106
rect 12014 31054 12066 31106
rect 12066 31054 12068 31106
rect 12012 31052 12068 31054
rect 12124 30940 12180 30996
rect 12684 53506 12740 53508
rect 12684 53454 12686 53506
rect 12686 53454 12738 53506
rect 12738 53454 12740 53506
rect 12684 53452 12740 53454
rect 12684 52108 12740 52164
rect 13804 53676 13860 53732
rect 12684 50482 12740 50484
rect 12684 50430 12686 50482
rect 12686 50430 12738 50482
rect 12738 50430 12740 50482
rect 12684 50428 12740 50430
rect 12796 48748 12852 48804
rect 12572 45948 12628 46004
rect 12684 43484 12740 43540
rect 12684 42588 12740 42644
rect 12684 38892 12740 38948
rect 13132 48636 13188 48692
rect 12908 43372 12964 43428
rect 12908 42700 12964 42756
rect 13804 48636 13860 48692
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 18732 55916 18788 55972
rect 18844 55804 18900 55860
rect 15260 55020 15316 55076
rect 14140 53058 14196 53060
rect 14140 53006 14142 53058
rect 14142 53006 14194 53058
rect 14194 53006 14196 53058
rect 14140 53004 14196 53006
rect 14812 53730 14868 53732
rect 14812 53678 14814 53730
rect 14814 53678 14866 53730
rect 14866 53678 14868 53730
rect 14812 53676 14868 53678
rect 15148 52220 15204 52276
rect 14476 52108 14532 52164
rect 15036 52108 15092 52164
rect 15036 49810 15092 49812
rect 15036 49758 15038 49810
rect 15038 49758 15090 49810
rect 15090 49758 15092 49810
rect 15036 49756 15092 49758
rect 16268 54460 16324 54516
rect 17948 55132 18004 55188
rect 17388 53676 17444 53732
rect 18732 55074 18788 55076
rect 18732 55022 18734 55074
rect 18734 55022 18786 55074
rect 18786 55022 18788 55074
rect 18732 55020 18788 55022
rect 18732 53730 18788 53732
rect 18732 53678 18734 53730
rect 18734 53678 18786 53730
rect 18786 53678 18788 53730
rect 18732 53676 18788 53678
rect 19292 54572 19348 54628
rect 28364 56140 28420 56196
rect 20636 55970 20692 55972
rect 20636 55918 20638 55970
rect 20638 55918 20690 55970
rect 20690 55918 20692 55970
rect 20636 55916 20692 55918
rect 22652 55804 22708 55860
rect 22764 55916 22820 55972
rect 18844 53564 18900 53620
rect 16492 52946 16548 52948
rect 16492 52894 16494 52946
rect 16494 52894 16546 52946
rect 16546 52894 16548 52946
rect 16492 52892 16548 52894
rect 16940 52220 16996 52276
rect 15820 52108 15876 52164
rect 16492 52162 16548 52164
rect 16492 52110 16494 52162
rect 16494 52110 16546 52162
rect 16546 52110 16548 52162
rect 16492 52108 16548 52110
rect 17052 52108 17108 52164
rect 17612 52108 17668 52164
rect 18172 52892 18228 52948
rect 15596 50594 15652 50596
rect 15596 50542 15598 50594
rect 15598 50542 15650 50594
rect 15650 50542 15652 50594
rect 15596 50540 15652 50542
rect 15260 49868 15316 49924
rect 15596 49756 15652 49812
rect 15596 48748 15652 48804
rect 15148 47964 15204 48020
rect 14028 47516 14084 47572
rect 16940 46508 16996 46564
rect 16156 45778 16212 45780
rect 16156 45726 16158 45778
rect 16158 45726 16210 45778
rect 16210 45726 16212 45778
rect 16156 45724 16212 45726
rect 14364 44098 14420 44100
rect 14364 44046 14366 44098
rect 14366 44046 14418 44098
rect 14418 44046 14420 44098
rect 14364 44044 14420 44046
rect 15372 44044 15428 44100
rect 16156 43762 16212 43764
rect 16156 43710 16158 43762
rect 16158 43710 16210 43762
rect 16210 43710 16212 43762
rect 16156 43708 16212 43710
rect 13580 43538 13636 43540
rect 13580 43486 13582 43538
rect 13582 43486 13634 43538
rect 13634 43486 13636 43538
rect 13580 43484 13636 43486
rect 13580 42754 13636 42756
rect 13580 42702 13582 42754
rect 13582 42702 13634 42754
rect 13634 42702 13636 42754
rect 13580 42700 13636 42702
rect 14252 42754 14308 42756
rect 14252 42702 14254 42754
rect 14254 42702 14306 42754
rect 14306 42702 14308 42754
rect 14252 42700 14308 42702
rect 15820 43148 15876 43204
rect 14924 41916 14980 41972
rect 15484 41132 15540 41188
rect 12796 37996 12852 38052
rect 13244 38892 13300 38948
rect 12908 37938 12964 37940
rect 12908 37886 12910 37938
rect 12910 37886 12962 37938
rect 12962 37886 12964 37938
rect 12908 37884 12964 37886
rect 12572 37266 12628 37268
rect 12572 37214 12574 37266
rect 12574 37214 12626 37266
rect 12626 37214 12628 37266
rect 12572 37212 12628 37214
rect 13692 38108 13748 38164
rect 14028 38108 14084 38164
rect 13356 37996 13412 38052
rect 13692 37884 13748 37940
rect 13132 37324 13188 37380
rect 12684 36876 12740 36932
rect 12460 36652 12516 36708
rect 13020 37154 13076 37156
rect 13020 37102 13022 37154
rect 13022 37102 13074 37154
rect 13074 37102 13076 37154
rect 13020 37100 13076 37102
rect 12796 36370 12852 36372
rect 12796 36318 12798 36370
rect 12798 36318 12850 36370
rect 12850 36318 12852 36370
rect 12796 36316 12852 36318
rect 12572 35868 12628 35924
rect 12460 35756 12516 35812
rect 12908 35810 12964 35812
rect 12908 35758 12910 35810
rect 12910 35758 12962 35810
rect 12962 35758 12964 35810
rect 12908 35756 12964 35758
rect 12572 35196 12628 35252
rect 12572 34748 12628 34804
rect 12460 32674 12516 32676
rect 12460 32622 12462 32674
rect 12462 32622 12514 32674
rect 12514 32622 12516 32674
rect 12460 32620 12516 32622
rect 13244 37100 13300 37156
rect 13468 36876 13524 36932
rect 12348 31554 12404 31556
rect 12348 31502 12350 31554
rect 12350 31502 12402 31554
rect 12402 31502 12404 31554
rect 12348 31500 12404 31502
rect 12348 30210 12404 30212
rect 12348 30158 12350 30210
rect 12350 30158 12402 30210
rect 12402 30158 12404 30210
rect 12348 30156 12404 30158
rect 12236 30098 12292 30100
rect 12236 30046 12238 30098
rect 12238 30046 12290 30098
rect 12290 30046 12292 30098
rect 12236 30044 12292 30046
rect 12236 29538 12292 29540
rect 12236 29486 12238 29538
rect 12238 29486 12290 29538
rect 12290 29486 12292 29538
rect 12236 29484 12292 29486
rect 12012 28588 12068 28644
rect 12348 28866 12404 28868
rect 12348 28814 12350 28866
rect 12350 28814 12402 28866
rect 12402 28814 12404 28866
rect 12348 28812 12404 28814
rect 12572 32396 12628 32452
rect 13244 36652 13300 36708
rect 13132 32450 13188 32452
rect 13132 32398 13134 32450
rect 13134 32398 13186 32450
rect 13186 32398 13188 32450
rect 13132 32396 13188 32398
rect 12684 31612 12740 31668
rect 12572 29932 12628 29988
rect 13020 31948 13076 32004
rect 13132 30156 13188 30212
rect 12796 30044 12852 30100
rect 12572 28754 12628 28756
rect 12572 28702 12574 28754
rect 12574 28702 12626 28754
rect 12626 28702 12628 28754
rect 12572 28700 12628 28702
rect 12460 28364 12516 28420
rect 11676 27074 11732 27076
rect 11676 27022 11678 27074
rect 11678 27022 11730 27074
rect 11730 27022 11732 27074
rect 11676 27020 11732 27022
rect 12124 27074 12180 27076
rect 12124 27022 12126 27074
rect 12126 27022 12178 27074
rect 12178 27022 12180 27074
rect 12124 27020 12180 27022
rect 14252 37884 14308 37940
rect 13468 36316 13524 36372
rect 13356 35586 13412 35588
rect 13356 35534 13358 35586
rect 13358 35534 13410 35586
rect 13410 35534 13412 35586
rect 13356 35532 13412 35534
rect 13580 32620 13636 32676
rect 16492 42642 16548 42644
rect 16492 42590 16494 42642
rect 16494 42590 16546 42642
rect 16546 42590 16548 42642
rect 16492 42588 16548 42590
rect 14588 37772 14644 37828
rect 14028 36876 14084 36932
rect 14140 36482 14196 36484
rect 14140 36430 14142 36482
rect 14142 36430 14194 36482
rect 14194 36430 14196 36482
rect 14140 36428 14196 36430
rect 15036 37100 15092 37156
rect 14476 35980 14532 36036
rect 15596 37826 15652 37828
rect 15596 37774 15598 37826
rect 15598 37774 15650 37826
rect 15650 37774 15652 37826
rect 15596 37772 15652 37774
rect 15372 37154 15428 37156
rect 15372 37102 15374 37154
rect 15374 37102 15426 37154
rect 15426 37102 15428 37154
rect 15372 37100 15428 37102
rect 15148 36428 15204 36484
rect 14140 35922 14196 35924
rect 14140 35870 14142 35922
rect 14142 35870 14194 35922
rect 14194 35870 14196 35922
rect 14140 35868 14196 35870
rect 14364 35868 14420 35924
rect 14700 35922 14756 35924
rect 14700 35870 14702 35922
rect 14702 35870 14754 35922
rect 14754 35870 14756 35922
rect 14700 35868 14756 35870
rect 14028 35532 14084 35588
rect 13916 31948 13972 32004
rect 13916 31612 13972 31668
rect 13244 29932 13300 29988
rect 13804 30098 13860 30100
rect 13804 30046 13806 30098
rect 13806 30046 13858 30098
rect 13858 30046 13860 30098
rect 13804 30044 13860 30046
rect 12908 28812 12964 28868
rect 15372 35810 15428 35812
rect 15372 35758 15374 35810
rect 15374 35758 15426 35810
rect 15426 35758 15428 35810
rect 15372 35756 15428 35758
rect 15148 35532 15204 35588
rect 15484 35644 15540 35700
rect 15820 35196 15876 35252
rect 16044 36258 16100 36260
rect 16044 36206 16046 36258
rect 16046 36206 16098 36258
rect 16098 36206 16100 36258
rect 16044 36204 16100 36206
rect 16044 35980 16100 36036
rect 16604 41916 16660 41972
rect 16716 41186 16772 41188
rect 16716 41134 16718 41186
rect 16718 41134 16770 41186
rect 16770 41134 16772 41186
rect 16716 41132 16772 41134
rect 16604 41020 16660 41076
rect 16604 40460 16660 40516
rect 16828 40796 16884 40852
rect 16492 38220 16548 38276
rect 17052 39004 17108 39060
rect 17164 39452 17220 39508
rect 16940 37490 16996 37492
rect 16940 37438 16942 37490
rect 16942 37438 16994 37490
rect 16994 37438 16996 37490
rect 16940 37436 16996 37438
rect 17388 41074 17444 41076
rect 17388 41022 17390 41074
rect 17390 41022 17442 41074
rect 17442 41022 17444 41074
rect 17388 41020 17444 41022
rect 17276 37996 17332 38052
rect 18060 51436 18116 51492
rect 18620 53058 18676 53060
rect 18620 53006 18622 53058
rect 18622 53006 18674 53058
rect 18674 53006 18676 53058
rect 18620 53004 18676 53006
rect 18284 52108 18340 52164
rect 18732 51490 18788 51492
rect 18732 51438 18734 51490
rect 18734 51438 18786 51490
rect 18786 51438 18788 51490
rect 18732 51436 18788 51438
rect 19404 54460 19460 54516
rect 18956 52220 19012 52276
rect 18620 50706 18676 50708
rect 18620 50654 18622 50706
rect 18622 50654 18674 50706
rect 18674 50654 18676 50706
rect 18620 50652 18676 50654
rect 18508 49756 18564 49812
rect 18172 48300 18228 48356
rect 18396 48748 18452 48804
rect 17724 44268 17780 44324
rect 17948 44156 18004 44212
rect 17724 43708 17780 43764
rect 17612 42754 17668 42756
rect 17612 42702 17614 42754
rect 17614 42702 17666 42754
rect 17666 42702 17668 42754
rect 17612 42700 17668 42702
rect 18060 42642 18116 42644
rect 18060 42590 18062 42642
rect 18062 42590 18114 42642
rect 18114 42590 18116 42642
rect 18060 42588 18116 42590
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 20188 54684 20244 54740
rect 20860 55074 20916 55076
rect 20860 55022 20862 55074
rect 20862 55022 20914 55074
rect 20914 55022 20916 55074
rect 20860 55020 20916 55022
rect 20300 54460 20356 54516
rect 19068 50204 19124 50260
rect 19180 50370 19236 50372
rect 19180 50318 19182 50370
rect 19182 50318 19234 50370
rect 19234 50318 19236 50370
rect 19180 50316 19236 50318
rect 18956 49810 19012 49812
rect 18956 49758 18958 49810
rect 18958 49758 19010 49810
rect 19010 49758 19012 49810
rect 18956 49756 19012 49758
rect 19180 49756 19236 49812
rect 20748 54348 20804 54404
rect 20860 53900 20916 53956
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19516 52780 19572 52836
rect 19964 52834 20020 52836
rect 19964 52782 19966 52834
rect 19966 52782 20018 52834
rect 20018 52782 20020 52834
rect 19964 52780 20020 52782
rect 20524 52780 20580 52836
rect 21532 52274 21588 52276
rect 21532 52222 21534 52274
rect 21534 52222 21586 52274
rect 21586 52222 21588 52274
rect 21532 52220 21588 52222
rect 21084 51996 21140 52052
rect 18844 44098 18900 44100
rect 18844 44046 18846 44098
rect 18846 44046 18898 44098
rect 18898 44046 18900 44098
rect 18844 44044 18900 44046
rect 18732 42476 18788 42532
rect 18620 40514 18676 40516
rect 18620 40462 18622 40514
rect 18622 40462 18674 40514
rect 18674 40462 18676 40514
rect 18620 40460 18676 40462
rect 17164 36876 17220 36932
rect 16492 36316 16548 36372
rect 16492 35756 16548 35812
rect 16268 35698 16324 35700
rect 16268 35646 16270 35698
rect 16270 35646 16322 35698
rect 16322 35646 16324 35698
rect 16268 35644 16324 35646
rect 16716 36204 16772 36260
rect 17388 36594 17444 36596
rect 17388 36542 17390 36594
rect 17390 36542 17442 36594
rect 17442 36542 17444 36594
rect 17388 36540 17444 36542
rect 16828 35644 16884 35700
rect 17724 37436 17780 37492
rect 17500 35868 17556 35924
rect 16044 35308 16100 35364
rect 16716 35420 16772 35476
rect 15820 34636 15876 34692
rect 16940 35308 16996 35364
rect 15148 32620 15204 32676
rect 16044 31890 16100 31892
rect 16044 31838 16046 31890
rect 16046 31838 16098 31890
rect 16098 31838 16100 31890
rect 16044 31836 16100 31838
rect 17276 35196 17332 35252
rect 17052 31836 17108 31892
rect 16604 31666 16660 31668
rect 16604 31614 16606 31666
rect 16606 31614 16658 31666
rect 16658 31614 16660 31666
rect 16604 31612 16660 31614
rect 17164 33404 17220 33460
rect 17724 36876 17780 36932
rect 17948 36652 18004 36708
rect 18172 37996 18228 38052
rect 17836 36428 17892 36484
rect 17836 36258 17892 36260
rect 17836 36206 17838 36258
rect 17838 36206 17890 36258
rect 17890 36206 17892 36258
rect 17836 36204 17892 36206
rect 17836 35644 17892 35700
rect 17836 35308 17892 35364
rect 17612 33404 17668 33460
rect 16044 31388 16100 31444
rect 16380 31388 16436 31444
rect 16044 30210 16100 30212
rect 16044 30158 16046 30210
rect 16046 30158 16098 30210
rect 16098 30158 16100 30210
rect 16044 30156 16100 30158
rect 14364 30044 14420 30100
rect 14924 30098 14980 30100
rect 14924 30046 14926 30098
rect 14926 30046 14978 30098
rect 14978 30046 14980 30098
rect 14924 30044 14980 30046
rect 15484 30098 15540 30100
rect 15484 30046 15486 30098
rect 15486 30046 15538 30098
rect 15538 30046 15540 30098
rect 15484 30044 15540 30046
rect 15484 29260 15540 29316
rect 13916 28812 13972 28868
rect 13580 28754 13636 28756
rect 13580 28702 13582 28754
rect 13582 28702 13634 28754
rect 13634 28702 13636 28754
rect 13580 28700 13636 28702
rect 17500 30492 17556 30548
rect 17052 30268 17108 30324
rect 16828 29820 16884 29876
rect 17164 30210 17220 30212
rect 17164 30158 17166 30210
rect 17166 30158 17218 30210
rect 17218 30158 17220 30210
rect 17164 30156 17220 30158
rect 16940 28754 16996 28756
rect 16940 28702 16942 28754
rect 16942 28702 16994 28754
rect 16994 28702 16996 28754
rect 16940 28700 16996 28702
rect 16604 28588 16660 28644
rect 17724 30322 17780 30324
rect 17724 30270 17726 30322
rect 17726 30270 17778 30322
rect 17778 30270 17780 30322
rect 17724 30268 17780 30270
rect 18060 36204 18116 36260
rect 18060 35308 18116 35364
rect 18284 36370 18340 36372
rect 18284 36318 18286 36370
rect 18286 36318 18338 36370
rect 18338 36318 18340 36370
rect 18284 36316 18340 36318
rect 18508 36988 18564 37044
rect 18284 35810 18340 35812
rect 18284 35758 18286 35810
rect 18286 35758 18338 35810
rect 18338 35758 18340 35810
rect 18284 35756 18340 35758
rect 18284 35308 18340 35364
rect 17948 30492 18004 30548
rect 18060 31612 18116 31668
rect 18060 30380 18116 30436
rect 17836 30156 17892 30212
rect 19516 50316 19572 50372
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19740 51548 19796 51604
rect 19740 50594 19796 50596
rect 19740 50542 19742 50594
rect 19742 50542 19794 50594
rect 19794 50542 19796 50594
rect 19740 50540 19796 50542
rect 20188 50316 20244 50372
rect 22092 50876 22148 50932
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19628 49644 19684 49700
rect 22652 52108 22708 52164
rect 24108 55804 24164 55860
rect 25340 56082 25396 56084
rect 25340 56030 25342 56082
rect 25342 56030 25394 56082
rect 25394 56030 25396 56082
rect 25340 56028 25396 56030
rect 24220 54402 24276 54404
rect 24220 54350 24222 54402
rect 24222 54350 24274 54402
rect 24274 54350 24276 54402
rect 24220 54348 24276 54350
rect 23212 53564 23268 53620
rect 23436 53170 23492 53172
rect 23436 53118 23438 53170
rect 23438 53118 23490 53170
rect 23490 53118 23492 53170
rect 23436 53116 23492 53118
rect 22204 49980 22260 50036
rect 20524 48748 20580 48804
rect 19404 47570 19460 47572
rect 19404 47518 19406 47570
rect 19406 47518 19458 47570
rect 19458 47518 19460 47570
rect 19404 47516 19460 47518
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19180 45890 19236 45892
rect 19180 45838 19182 45890
rect 19182 45838 19234 45890
rect 19234 45838 19236 45890
rect 19180 45836 19236 45838
rect 19404 45612 19460 45668
rect 19292 44210 19348 44212
rect 19292 44158 19294 44210
rect 19294 44158 19346 44210
rect 19346 44158 19348 44210
rect 19292 44156 19348 44158
rect 18956 40908 19012 40964
rect 19068 40460 19124 40516
rect 18956 37436 19012 37492
rect 18844 37212 18900 37268
rect 18732 36988 18788 37044
rect 18732 36204 18788 36260
rect 18508 34802 18564 34804
rect 18508 34750 18510 34802
rect 18510 34750 18562 34802
rect 18562 34750 18564 34802
rect 18508 34748 18564 34750
rect 18620 33180 18676 33236
rect 18620 30210 18676 30212
rect 18620 30158 18622 30210
rect 18622 30158 18674 30210
rect 18674 30158 18676 30210
rect 18620 30156 18676 30158
rect 18284 29820 18340 29876
rect 18508 29986 18564 29988
rect 18508 29934 18510 29986
rect 18510 29934 18562 29986
rect 18562 29934 18564 29986
rect 18508 29932 18564 29934
rect 19292 37436 19348 37492
rect 20076 46562 20132 46564
rect 20076 46510 20078 46562
rect 20078 46510 20130 46562
rect 20130 46510 20132 46562
rect 20076 46508 20132 46510
rect 19740 45612 19796 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19628 44044 19684 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 21532 48802 21588 48804
rect 21532 48750 21534 48802
rect 21534 48750 21586 48802
rect 21586 48750 21588 48802
rect 21532 48748 21588 48750
rect 22204 48748 22260 48804
rect 23100 49698 23156 49700
rect 23100 49646 23102 49698
rect 23102 49646 23154 49698
rect 23154 49646 23156 49698
rect 23100 49644 23156 49646
rect 21084 46396 21140 46452
rect 21868 45948 21924 46004
rect 20860 45836 20916 45892
rect 20748 45106 20804 45108
rect 20748 45054 20750 45106
rect 20750 45054 20802 45106
rect 20802 45054 20804 45106
rect 20748 45052 20804 45054
rect 20524 41132 20580 41188
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19628 40460 19684 40516
rect 20636 40460 20692 40516
rect 19516 39564 19572 39620
rect 19740 40236 19796 40292
rect 20076 39842 20132 39844
rect 20076 39790 20078 39842
rect 20078 39790 20130 39842
rect 20130 39790 20132 39842
rect 20076 39788 20132 39790
rect 20748 40124 20804 40180
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20412 39058 20468 39060
rect 20412 39006 20414 39058
rect 20414 39006 20466 39058
rect 20466 39006 20468 39058
rect 20412 39004 20468 39006
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20524 37490 20580 37492
rect 20524 37438 20526 37490
rect 20526 37438 20578 37490
rect 20578 37438 20580 37490
rect 20524 37436 20580 37438
rect 19068 36594 19124 36596
rect 19068 36542 19070 36594
rect 19070 36542 19122 36594
rect 19122 36542 19124 36594
rect 19068 36540 19124 36542
rect 19180 36482 19236 36484
rect 19180 36430 19182 36482
rect 19182 36430 19234 36482
rect 19234 36430 19236 36482
rect 19180 36428 19236 36430
rect 18956 36258 19012 36260
rect 18956 36206 18958 36258
rect 18958 36206 19010 36258
rect 19010 36206 19012 36258
rect 18956 36204 19012 36206
rect 19180 36092 19236 36148
rect 19068 34802 19124 34804
rect 19068 34750 19070 34802
rect 19070 34750 19122 34802
rect 19122 34750 19124 34802
rect 19068 34748 19124 34750
rect 18844 33292 18900 33348
rect 19740 37266 19796 37268
rect 19740 37214 19742 37266
rect 19742 37214 19794 37266
rect 19794 37214 19796 37266
rect 19740 37212 19796 37214
rect 19964 36988 20020 37044
rect 19404 36482 19460 36484
rect 19404 36430 19406 36482
rect 19406 36430 19458 36482
rect 19458 36430 19460 36482
rect 19404 36428 19460 36430
rect 19852 36594 19908 36596
rect 19852 36542 19854 36594
rect 19854 36542 19906 36594
rect 19906 36542 19908 36594
rect 19852 36540 19908 36542
rect 20412 36594 20468 36596
rect 20412 36542 20414 36594
rect 20414 36542 20466 36594
rect 20466 36542 20468 36594
rect 20412 36540 20468 36542
rect 19292 35868 19348 35924
rect 19292 35698 19348 35700
rect 19292 35646 19294 35698
rect 19294 35646 19346 35698
rect 19346 35646 19348 35698
rect 19292 35644 19348 35646
rect 19516 35308 19572 35364
rect 20188 36204 20244 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20076 35922 20132 35924
rect 20076 35870 20078 35922
rect 20078 35870 20130 35922
rect 20130 35870 20132 35922
rect 20076 35868 20132 35870
rect 19852 35756 19908 35812
rect 20972 43596 21028 43652
rect 21532 41186 21588 41188
rect 21532 41134 21534 41186
rect 21534 41134 21586 41186
rect 21586 41134 21588 41186
rect 21532 41132 21588 41134
rect 21532 39618 21588 39620
rect 21532 39566 21534 39618
rect 21534 39566 21586 39618
rect 21586 39566 21588 39618
rect 21532 39564 21588 39566
rect 21756 39004 21812 39060
rect 20972 37266 21028 37268
rect 20972 37214 20974 37266
rect 20974 37214 21026 37266
rect 21026 37214 21028 37266
rect 20972 37212 21028 37214
rect 21756 35868 21812 35924
rect 19292 34690 19348 34692
rect 19292 34638 19294 34690
rect 19294 34638 19346 34690
rect 19346 34638 19348 34690
rect 19292 34636 19348 34638
rect 19852 34690 19908 34692
rect 19852 34638 19854 34690
rect 19854 34638 19906 34690
rect 19906 34638 19908 34690
rect 19852 34636 19908 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19404 33964 19460 34020
rect 19852 34018 19908 34020
rect 19852 33966 19854 34018
rect 19854 33966 19906 34018
rect 19906 33966 19908 34018
rect 19852 33964 19908 33966
rect 19964 33906 20020 33908
rect 19964 33854 19966 33906
rect 19966 33854 20018 33906
rect 20018 33854 20020 33906
rect 19964 33852 20020 33854
rect 20412 34860 20468 34916
rect 20188 33852 20244 33908
rect 20860 34690 20916 34692
rect 20860 34638 20862 34690
rect 20862 34638 20914 34690
rect 20914 34638 20916 34690
rect 20860 34636 20916 34638
rect 20524 34188 20580 34244
rect 20412 34018 20468 34020
rect 20412 33966 20414 34018
rect 20414 33966 20466 34018
rect 20466 33966 20468 34018
rect 20412 33964 20468 33966
rect 20300 33628 20356 33684
rect 19292 33068 19348 33124
rect 18396 29596 18452 29652
rect 18956 30044 19012 30100
rect 18284 29538 18340 29540
rect 18284 29486 18286 29538
rect 18286 29486 18338 29538
rect 18338 29486 18340 29538
rect 18284 29484 18340 29486
rect 17948 28812 18004 28868
rect 18172 28642 18228 28644
rect 18172 28590 18174 28642
rect 18174 28590 18226 28642
rect 18226 28590 18228 28642
rect 18172 28588 18228 28590
rect 17724 28476 17780 28532
rect 18508 28700 18564 28756
rect 17388 27074 17444 27076
rect 17388 27022 17390 27074
rect 17390 27022 17442 27074
rect 17442 27022 17444 27074
rect 17388 27020 17444 27022
rect 11340 26572 11396 26628
rect 18284 27186 18340 27188
rect 18284 27134 18286 27186
rect 18286 27134 18338 27186
rect 18338 27134 18340 27186
rect 18284 27132 18340 27134
rect 17836 26908 17892 26964
rect 12012 26684 12068 26740
rect 11900 26066 11956 26068
rect 11900 26014 11902 26066
rect 11902 26014 11954 26066
rect 11954 26014 11956 26066
rect 11900 26012 11956 26014
rect 11340 24834 11396 24836
rect 11340 24782 11342 24834
rect 11342 24782 11394 24834
rect 11394 24782 11396 24834
rect 11340 24780 11396 24782
rect 11116 24722 11172 24724
rect 11116 24670 11118 24722
rect 11118 24670 11170 24722
rect 11170 24670 11172 24722
rect 11116 24668 11172 24670
rect 11788 24668 11844 24724
rect 11340 23436 11396 23492
rect 10668 23042 10724 23044
rect 10668 22990 10670 23042
rect 10670 22990 10722 23042
rect 10722 22990 10724 23042
rect 10668 22988 10724 22990
rect 11004 22988 11060 23044
rect 11676 23042 11732 23044
rect 11676 22990 11678 23042
rect 11678 22990 11730 23042
rect 11730 22990 11732 23042
rect 11676 22988 11732 22990
rect 12236 24834 12292 24836
rect 12236 24782 12238 24834
rect 12238 24782 12290 24834
rect 12290 24782 12292 24834
rect 12236 24780 12292 24782
rect 9996 22258 10052 22260
rect 9996 22206 9998 22258
rect 9998 22206 10050 22258
rect 10050 22206 10052 22258
rect 9996 22204 10052 22206
rect 9436 21756 9492 21812
rect 11676 22316 11732 22372
rect 7532 12348 7588 12404
rect 6412 6076 6468 6132
rect 11340 5292 11396 5348
rect 12236 22370 12292 22372
rect 12236 22318 12238 22370
rect 12238 22318 12290 22370
rect 12290 22318 12292 22370
rect 12236 22316 12292 22318
rect 11788 22204 11844 22260
rect 11116 4562 11172 4564
rect 11116 4510 11118 4562
rect 11118 4510 11170 4562
rect 11170 4510 11172 4562
rect 11116 4508 11172 4510
rect 12460 26684 12516 26740
rect 18172 24780 18228 24836
rect 18060 24556 18116 24612
rect 17164 23436 17220 23492
rect 17724 23826 17780 23828
rect 17724 23774 17726 23826
rect 17726 23774 17778 23826
rect 17778 23774 17780 23826
rect 17724 23772 17780 23774
rect 17948 23436 18004 23492
rect 17388 23324 17444 23380
rect 17836 23324 17892 23380
rect 19180 30434 19236 30436
rect 19180 30382 19182 30434
rect 19182 30382 19234 30434
rect 19234 30382 19236 30434
rect 19180 30380 19236 30382
rect 19068 29596 19124 29652
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19628 30210 19684 30212
rect 19628 30158 19630 30210
rect 19630 30158 19682 30210
rect 19682 30158 19684 30210
rect 19628 30156 19684 30158
rect 19964 30098 20020 30100
rect 19964 30046 19966 30098
rect 19966 30046 20018 30098
rect 20018 30046 20020 30098
rect 19964 30044 20020 30046
rect 20412 30044 20468 30100
rect 20412 29820 20468 29876
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18732 28700 18788 28756
rect 19516 29538 19572 29540
rect 19516 29486 19518 29538
rect 19518 29486 19570 29538
rect 19570 29486 19572 29538
rect 19516 29484 19572 29486
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 27804 19572 27860
rect 19180 27132 19236 27188
rect 19404 27132 19460 27188
rect 20188 27692 20244 27748
rect 22204 40626 22260 40628
rect 22204 40574 22206 40626
rect 22206 40574 22258 40626
rect 22258 40574 22260 40626
rect 22204 40572 22260 40574
rect 23660 50316 23716 50372
rect 23660 49756 23716 49812
rect 23212 48076 23268 48132
rect 23436 47180 23492 47236
rect 23324 47068 23380 47124
rect 23548 46396 23604 46452
rect 23436 43762 23492 43764
rect 23436 43710 23438 43762
rect 23438 43710 23490 43762
rect 23490 43710 23492 43762
rect 23436 43708 23492 43710
rect 23212 42194 23268 42196
rect 23212 42142 23214 42194
rect 23214 42142 23266 42194
rect 23266 42142 23268 42194
rect 23212 42140 23268 42142
rect 22764 41132 22820 41188
rect 23212 40236 23268 40292
rect 23212 38780 23268 38836
rect 22540 35196 22596 35252
rect 22428 35026 22484 35028
rect 22428 34974 22430 35026
rect 22430 34974 22482 35026
rect 22482 34974 22484 35026
rect 22428 34972 22484 34974
rect 22092 34914 22148 34916
rect 22092 34862 22094 34914
rect 22094 34862 22146 34914
rect 22146 34862 22148 34914
rect 22092 34860 22148 34862
rect 21756 34524 21812 34580
rect 21980 34690 22036 34692
rect 21980 34638 21982 34690
rect 21982 34638 22034 34690
rect 22034 34638 22036 34690
rect 21980 34636 22036 34638
rect 21644 33852 21700 33908
rect 21420 32562 21476 32564
rect 21420 32510 21422 32562
rect 21422 32510 21474 32562
rect 21474 32510 21476 32562
rect 21420 32508 21476 32510
rect 20972 31724 21028 31780
rect 21644 30210 21700 30212
rect 21644 30158 21646 30210
rect 21646 30158 21698 30210
rect 21698 30158 21700 30210
rect 21644 30156 21700 30158
rect 20860 30098 20916 30100
rect 20860 30046 20862 30098
rect 20862 30046 20914 30098
rect 20914 30046 20916 30098
rect 20860 30044 20916 30046
rect 20860 29484 20916 29540
rect 21868 29820 21924 29876
rect 20524 27692 20580 27748
rect 22316 33292 22372 33348
rect 22204 32562 22260 32564
rect 22204 32510 22206 32562
rect 22206 32510 22258 32562
rect 22258 32510 22260 32562
rect 22204 32508 22260 32510
rect 22092 29932 22148 29988
rect 22652 32396 22708 32452
rect 23100 37772 23156 37828
rect 22876 36258 22932 36260
rect 22876 36206 22878 36258
rect 22878 36206 22930 36258
rect 22930 36206 22932 36258
rect 22876 36204 22932 36206
rect 22988 35026 23044 35028
rect 22988 34974 22990 35026
rect 22990 34974 23042 35026
rect 23042 34974 23044 35026
rect 22988 34972 23044 34974
rect 24108 52722 24164 52724
rect 24108 52670 24110 52722
rect 24110 52670 24162 52722
rect 24162 52670 24164 52722
rect 24108 52668 24164 52670
rect 26796 56082 26852 56084
rect 26796 56030 26798 56082
rect 26798 56030 26850 56082
rect 26850 56030 26852 56082
rect 26796 56028 26852 56030
rect 27356 53618 27412 53620
rect 27356 53566 27358 53618
rect 27358 53566 27410 53618
rect 27410 53566 27412 53618
rect 27356 53564 27412 53566
rect 27804 53564 27860 53620
rect 27356 52834 27412 52836
rect 27356 52782 27358 52834
rect 27358 52782 27410 52834
rect 27410 52782 27412 52834
rect 27356 52780 27412 52782
rect 25340 52668 25396 52724
rect 25900 52668 25956 52724
rect 24556 51996 24612 52052
rect 25228 51996 25284 52052
rect 24556 46396 24612 46452
rect 24108 46284 24164 46340
rect 23660 40626 23716 40628
rect 23660 40574 23662 40626
rect 23662 40574 23714 40626
rect 23714 40574 23716 40626
rect 23660 40572 23716 40574
rect 23772 39116 23828 39172
rect 23548 36876 23604 36932
rect 22876 32284 22932 32340
rect 22764 30044 22820 30100
rect 22316 29820 22372 29876
rect 22092 29708 22148 29764
rect 22204 29596 22260 29652
rect 21980 27580 22036 27636
rect 20188 27186 20244 27188
rect 20188 27134 20190 27186
rect 20190 27134 20242 27186
rect 20242 27134 20244 27186
rect 20188 27132 20244 27134
rect 19628 27074 19684 27076
rect 19628 27022 19630 27074
rect 19630 27022 19682 27074
rect 19682 27022 19684 27074
rect 21868 27132 21924 27188
rect 19628 27020 19684 27022
rect 19516 26962 19572 26964
rect 19516 26910 19518 26962
rect 19518 26910 19570 26962
rect 19570 26910 19572 26962
rect 19516 26908 19572 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 25228 19684 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19628 24610 19684 24612
rect 19628 24558 19630 24610
rect 19630 24558 19682 24610
rect 19682 24558 19684 24610
rect 19628 24556 19684 24558
rect 21868 24556 21924 24612
rect 21196 23660 21252 23716
rect 19836 23546 19892 23548
rect 18620 23436 18676 23492
rect 19180 23436 19236 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18172 23324 18228 23380
rect 18844 23378 18900 23380
rect 18844 23326 18846 23378
rect 18846 23326 18898 23378
rect 18898 23326 18900 23378
rect 18844 23324 18900 23326
rect 21644 23714 21700 23716
rect 21644 23662 21646 23714
rect 21646 23662 21698 23714
rect 21698 23662 21700 23714
rect 21644 23660 21700 23662
rect 16940 23042 16996 23044
rect 16940 22990 16942 23042
rect 16942 22990 16994 23042
rect 16994 22990 16996 23042
rect 16940 22988 16996 22990
rect 18396 22988 18452 23044
rect 21644 23042 21700 23044
rect 21644 22990 21646 23042
rect 21646 22990 21698 23042
rect 21698 22990 21700 23042
rect 21644 22988 21700 22990
rect 23548 36204 23604 36260
rect 23324 34524 23380 34580
rect 23324 32284 23380 32340
rect 23772 34188 23828 34244
rect 23996 43314 24052 43316
rect 23996 43262 23998 43314
rect 23998 43262 24050 43314
rect 24050 43262 24052 43314
rect 23996 43260 24052 43262
rect 24892 45164 24948 45220
rect 24332 45052 24388 45108
rect 24332 43650 24388 43652
rect 24332 43598 24334 43650
rect 24334 43598 24386 43650
rect 24386 43598 24388 43650
rect 24332 43596 24388 43598
rect 24220 40124 24276 40180
rect 24332 40908 24388 40964
rect 24108 40012 24164 40068
rect 24108 37996 24164 38052
rect 24108 37324 24164 37380
rect 24108 36370 24164 36372
rect 24108 36318 24110 36370
rect 24110 36318 24162 36370
rect 24162 36318 24164 36370
rect 24108 36316 24164 36318
rect 24220 34690 24276 34692
rect 24220 34638 24222 34690
rect 24222 34638 24274 34690
rect 24274 34638 24276 34690
rect 24220 34636 24276 34638
rect 23884 34076 23940 34132
rect 23996 33458 24052 33460
rect 23996 33406 23998 33458
rect 23998 33406 24050 33458
rect 24050 33406 24052 33458
rect 23996 33404 24052 33406
rect 24892 43708 24948 43764
rect 24668 42140 24724 42196
rect 24556 38162 24612 38164
rect 24556 38110 24558 38162
rect 24558 38110 24610 38162
rect 24610 38110 24612 38162
rect 24556 38108 24612 38110
rect 24444 36876 24500 36932
rect 25004 37826 25060 37828
rect 25004 37774 25006 37826
rect 25006 37774 25058 37826
rect 25058 37774 25060 37826
rect 25004 37772 25060 37774
rect 25004 37378 25060 37380
rect 25004 37326 25006 37378
rect 25006 37326 25058 37378
rect 25058 37326 25060 37378
rect 25004 37324 25060 37326
rect 25116 36428 25172 36484
rect 24892 36316 24948 36372
rect 24780 36258 24836 36260
rect 24780 36206 24782 36258
rect 24782 36206 24834 36258
rect 24834 36206 24836 36258
rect 24780 36204 24836 36206
rect 24892 35420 24948 35476
rect 25004 35084 25060 35140
rect 25004 34914 25060 34916
rect 25004 34862 25006 34914
rect 25006 34862 25058 34914
rect 25058 34862 25060 34914
rect 25004 34860 25060 34862
rect 25228 36316 25284 36372
rect 27244 50876 27300 50932
rect 26572 48188 26628 48244
rect 26348 40684 26404 40740
rect 25900 40460 25956 40516
rect 26012 39340 26068 39396
rect 25676 38108 25732 38164
rect 25564 38050 25620 38052
rect 25564 37998 25566 38050
rect 25566 37998 25618 38050
rect 25618 37998 25620 38050
rect 25564 37996 25620 37998
rect 25900 37938 25956 37940
rect 25900 37886 25902 37938
rect 25902 37886 25954 37938
rect 25954 37886 25956 37938
rect 25900 37884 25956 37886
rect 26124 38050 26180 38052
rect 26124 37998 26126 38050
rect 26126 37998 26178 38050
rect 26178 37998 26180 38050
rect 26124 37996 26180 37998
rect 26124 37772 26180 37828
rect 25788 37378 25844 37380
rect 25788 37326 25790 37378
rect 25790 37326 25842 37378
rect 25842 37326 25844 37378
rect 25788 37324 25844 37326
rect 25676 37266 25732 37268
rect 25676 37214 25678 37266
rect 25678 37214 25730 37266
rect 25730 37214 25732 37266
rect 26348 39394 26404 39396
rect 26348 39342 26350 39394
rect 26350 39342 26402 39394
rect 26402 39342 26404 39394
rect 26348 39340 26404 39342
rect 25676 37212 25732 37214
rect 25676 36988 25732 37044
rect 26460 38444 26516 38500
rect 25676 35980 25732 36036
rect 25452 35308 25508 35364
rect 26236 35980 26292 36036
rect 26012 35532 26068 35588
rect 24444 33292 24500 33348
rect 23772 32450 23828 32452
rect 23772 32398 23774 32450
rect 23774 32398 23826 32450
rect 23826 32398 23828 32450
rect 23772 32396 23828 32398
rect 24108 32284 24164 32340
rect 23884 31500 23940 31556
rect 23660 31164 23716 31220
rect 23548 29484 23604 29540
rect 23100 29036 23156 29092
rect 23100 28642 23156 28644
rect 23100 28590 23102 28642
rect 23102 28590 23154 28642
rect 23154 28590 23156 28642
rect 23100 28588 23156 28590
rect 22316 27244 22372 27300
rect 22428 28028 22484 28084
rect 23436 29036 23492 29092
rect 23324 28812 23380 28868
rect 23436 28642 23492 28644
rect 23436 28590 23438 28642
rect 23438 28590 23490 28642
rect 23490 28590 23492 28642
rect 23436 28588 23492 28590
rect 23548 28476 23604 28532
rect 23772 27970 23828 27972
rect 23772 27918 23774 27970
rect 23774 27918 23826 27970
rect 23826 27918 23828 27970
rect 23772 27916 23828 27918
rect 23548 27580 23604 27636
rect 22428 27132 22484 27188
rect 23324 27468 23380 27524
rect 22540 26908 22596 26964
rect 22428 25618 22484 25620
rect 22428 25566 22430 25618
rect 22430 25566 22482 25618
rect 22482 25566 22484 25618
rect 22428 25564 22484 25566
rect 23212 27020 23268 27076
rect 23436 27356 23492 27412
rect 24332 31554 24388 31556
rect 24332 31502 24334 31554
rect 24334 31502 24386 31554
rect 24386 31502 24388 31554
rect 24332 31500 24388 31502
rect 24220 28812 24276 28868
rect 24220 28476 24276 28532
rect 24108 27916 24164 27972
rect 22988 25618 23044 25620
rect 22988 25566 22990 25618
rect 22990 25566 23042 25618
rect 23042 25566 23044 25618
rect 22988 25564 23044 25566
rect 22876 25228 22932 25284
rect 23996 27468 24052 27524
rect 24444 27132 24500 27188
rect 25452 34802 25508 34804
rect 25452 34750 25454 34802
rect 25454 34750 25506 34802
rect 25506 34750 25508 34802
rect 25452 34748 25508 34750
rect 25228 34636 25284 34692
rect 25116 34076 25172 34132
rect 25004 33122 25060 33124
rect 25004 33070 25006 33122
rect 25006 33070 25058 33122
rect 25058 33070 25060 33122
rect 25004 33068 25060 33070
rect 25004 32508 25060 32564
rect 24780 31164 24836 31220
rect 24668 28642 24724 28644
rect 24668 28590 24670 28642
rect 24670 28590 24722 28642
rect 24722 28590 24724 28642
rect 24668 28588 24724 28590
rect 24668 27580 24724 27636
rect 24892 29650 24948 29652
rect 24892 29598 24894 29650
rect 24894 29598 24946 29650
rect 24946 29598 24948 29650
rect 24892 29596 24948 29598
rect 24668 26962 24724 26964
rect 24668 26910 24670 26962
rect 24670 26910 24722 26962
rect 24722 26910 24724 26962
rect 24668 26908 24724 26910
rect 25228 33628 25284 33684
rect 25676 34188 25732 34244
rect 25452 33458 25508 33460
rect 25452 33406 25454 33458
rect 25454 33406 25506 33458
rect 25506 33406 25508 33458
rect 25452 33404 25508 33406
rect 25564 33068 25620 33124
rect 26236 35308 26292 35364
rect 26012 33404 26068 33460
rect 26124 33964 26180 34020
rect 25788 33346 25844 33348
rect 25788 33294 25790 33346
rect 25790 33294 25842 33346
rect 25842 33294 25844 33346
rect 25788 33292 25844 33294
rect 25676 32620 25732 32676
rect 26012 32284 26068 32340
rect 25340 30828 25396 30884
rect 25116 27356 25172 27412
rect 25228 28588 25284 28644
rect 25116 27074 25172 27076
rect 25116 27022 25118 27074
rect 25118 27022 25170 27074
rect 25170 27022 25172 27074
rect 25116 27020 25172 27022
rect 26348 34914 26404 34916
rect 26348 34862 26350 34914
rect 26350 34862 26402 34914
rect 26402 34862 26404 34914
rect 26348 34860 26404 34862
rect 26348 34188 26404 34244
rect 26796 47570 26852 47572
rect 26796 47518 26798 47570
rect 26798 47518 26850 47570
rect 26850 47518 26852 47570
rect 26796 47516 26852 47518
rect 28028 53058 28084 53060
rect 28028 53006 28030 53058
rect 28030 53006 28082 53058
rect 28082 53006 28084 53058
rect 28028 53004 28084 53006
rect 28588 55132 28644 55188
rect 31836 56194 31892 56196
rect 31836 56142 31838 56194
rect 31838 56142 31890 56194
rect 31890 56142 31892 56194
rect 31836 56140 31892 56142
rect 31500 56028 31556 56084
rect 32060 56082 32116 56084
rect 32060 56030 32062 56082
rect 32062 56030 32114 56082
rect 32114 56030 32116 56082
rect 32060 56028 32116 56030
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 38220 56194 38276 56196
rect 38220 56142 38222 56194
rect 38222 56142 38274 56194
rect 38274 56142 38276 56194
rect 38220 56140 38276 56142
rect 39788 56140 39844 56196
rect 29260 55132 29316 55188
rect 28476 54572 28532 54628
rect 27356 47570 27412 47572
rect 27356 47518 27358 47570
rect 27358 47518 27410 47570
rect 27410 47518 27412 47570
rect 27356 47516 27412 47518
rect 28700 54236 28756 54292
rect 28812 53618 28868 53620
rect 28812 53566 28814 53618
rect 28814 53566 28866 53618
rect 28866 53566 28868 53618
rect 28812 53564 28868 53566
rect 30268 53954 30324 53956
rect 30268 53902 30270 53954
rect 30270 53902 30322 53954
rect 30322 53902 30324 53954
rect 30268 53900 30324 53902
rect 29148 53564 29204 53620
rect 29484 53564 29540 53620
rect 30380 53618 30436 53620
rect 30380 53566 30382 53618
rect 30382 53566 30434 53618
rect 30434 53566 30436 53618
rect 30380 53564 30436 53566
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 32508 53730 32564 53732
rect 32508 53678 32510 53730
rect 32510 53678 32562 53730
rect 32562 53678 32564 53730
rect 32508 53676 32564 53678
rect 30716 53564 30772 53620
rect 31052 53618 31108 53620
rect 31052 53566 31054 53618
rect 31054 53566 31106 53618
rect 31106 53566 31108 53618
rect 31052 53564 31108 53566
rect 29036 53170 29092 53172
rect 29036 53118 29038 53170
rect 29038 53118 29090 53170
rect 29090 53118 29092 53170
rect 29036 53116 29092 53118
rect 27916 47234 27972 47236
rect 27916 47182 27918 47234
rect 27918 47182 27970 47234
rect 27970 47182 27972 47234
rect 27916 47180 27972 47182
rect 28476 52274 28532 52276
rect 28476 52222 28478 52274
rect 28478 52222 28530 52274
rect 28530 52222 28532 52274
rect 28476 52220 28532 52222
rect 29148 52220 29204 52276
rect 30492 53452 30548 53508
rect 29708 53228 29764 53284
rect 29484 52274 29540 52276
rect 29484 52222 29486 52274
rect 29486 52222 29538 52274
rect 29538 52222 29540 52274
rect 29484 52220 29540 52222
rect 29820 52834 29876 52836
rect 29820 52782 29822 52834
rect 29822 52782 29874 52834
rect 29874 52782 29876 52834
rect 29820 52780 29876 52782
rect 30044 52274 30100 52276
rect 30044 52222 30046 52274
rect 30046 52222 30098 52274
rect 30098 52222 30100 52274
rect 30044 52220 30100 52222
rect 28364 52162 28420 52164
rect 28364 52110 28366 52162
rect 28366 52110 28418 52162
rect 28418 52110 28420 52162
rect 28364 52108 28420 52110
rect 30940 52892 30996 52948
rect 30716 52108 30772 52164
rect 31388 52556 31444 52612
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 32620 52220 32676 52276
rect 31052 51436 31108 51492
rect 30380 51324 30436 51380
rect 29820 51100 29876 51156
rect 28028 46956 28084 47012
rect 28364 49644 28420 49700
rect 27580 45330 27636 45332
rect 27580 45278 27582 45330
rect 27582 45278 27634 45330
rect 27634 45278 27636 45330
rect 27580 45276 27636 45278
rect 27244 42140 27300 42196
rect 26796 41020 26852 41076
rect 27244 40460 27300 40516
rect 26908 40236 26964 40292
rect 27468 40514 27524 40516
rect 27468 40462 27470 40514
rect 27470 40462 27522 40514
rect 27522 40462 27524 40514
rect 27468 40460 27524 40462
rect 27356 40290 27412 40292
rect 27356 40238 27358 40290
rect 27358 40238 27410 40290
rect 27410 40238 27412 40290
rect 27356 40236 27412 40238
rect 27916 44994 27972 44996
rect 27916 44942 27918 44994
rect 27918 44942 27970 44994
rect 27970 44942 27972 44994
rect 27916 44940 27972 44942
rect 27916 41020 27972 41076
rect 27692 40572 27748 40628
rect 27804 40684 27860 40740
rect 27916 40572 27972 40628
rect 28252 46956 28308 47012
rect 29596 48748 29652 48804
rect 28588 47068 28644 47124
rect 28700 46956 28756 47012
rect 29484 46956 29540 47012
rect 29372 46562 29428 46564
rect 29372 46510 29374 46562
rect 29374 46510 29426 46562
rect 29426 46510 29428 46562
rect 29372 46508 29428 46510
rect 28588 45164 28644 45220
rect 28700 45052 28756 45108
rect 29260 45276 29316 45332
rect 28140 40236 28196 40292
rect 26796 39394 26852 39396
rect 26796 39342 26798 39394
rect 26798 39342 26850 39394
rect 26850 39342 26852 39394
rect 26796 39340 26852 39342
rect 28812 44434 28868 44436
rect 28812 44382 28814 44434
rect 28814 44382 28866 44434
rect 28866 44382 28868 44434
rect 28812 44380 28868 44382
rect 28476 42588 28532 42644
rect 29596 44492 29652 44548
rect 29708 45106 29764 45108
rect 29708 45054 29710 45106
rect 29710 45054 29762 45106
rect 29762 45054 29764 45106
rect 29708 45052 29764 45054
rect 29484 42140 29540 42196
rect 28364 41244 28420 41300
rect 28812 41298 28868 41300
rect 28812 41246 28814 41298
rect 28814 41246 28866 41298
rect 28866 41246 28868 41298
rect 28812 41244 28868 41246
rect 29708 41132 29764 41188
rect 30380 49868 30436 49924
rect 32172 49922 32228 49924
rect 32172 49870 32174 49922
rect 32174 49870 32226 49922
rect 32226 49870 32228 49922
rect 32172 49868 32228 49870
rect 29932 46956 29988 47012
rect 29932 45330 29988 45332
rect 29932 45278 29934 45330
rect 29934 45278 29986 45330
rect 29986 45278 29988 45330
rect 29932 45276 29988 45278
rect 30268 45164 30324 45220
rect 29820 41244 29876 41300
rect 29932 44940 29988 44996
rect 30156 44940 30212 44996
rect 30156 44546 30212 44548
rect 30156 44494 30158 44546
rect 30158 44494 30210 44546
rect 30210 44494 30212 44546
rect 30156 44492 30212 44494
rect 31500 49698 31556 49700
rect 31500 49646 31502 49698
rect 31502 49646 31554 49698
rect 31554 49646 31556 49698
rect 31500 49644 31556 49646
rect 31388 48412 31444 48468
rect 32396 49868 32452 49924
rect 32172 49644 32228 49700
rect 32060 49586 32116 49588
rect 32060 49534 32062 49586
rect 32062 49534 32114 49586
rect 32114 49534 32116 49586
rect 32060 49532 32116 49534
rect 35532 52108 35588 52164
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 32620 49922 32676 49924
rect 32620 49870 32622 49922
rect 32622 49870 32674 49922
rect 32674 49870 32676 49922
rect 32620 49868 32676 49870
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 32508 49084 32564 49140
rect 31836 48914 31892 48916
rect 31836 48862 31838 48914
rect 31838 48862 31890 48914
rect 31890 48862 31892 48914
rect 31836 48860 31892 48862
rect 31612 47404 31668 47460
rect 30716 45890 30772 45892
rect 30716 45838 30718 45890
rect 30718 45838 30770 45890
rect 30770 45838 30772 45890
rect 30716 45836 30772 45838
rect 31164 45836 31220 45892
rect 30380 45052 30436 45108
rect 30268 44434 30324 44436
rect 30268 44382 30270 44434
rect 30270 44382 30322 44434
rect 30322 44382 30324 44434
rect 30268 44380 30324 44382
rect 30044 43596 30100 43652
rect 30940 45388 30996 45444
rect 30716 45330 30772 45332
rect 30716 45278 30718 45330
rect 30718 45278 30770 45330
rect 30770 45278 30772 45330
rect 30716 45276 30772 45278
rect 30604 45164 30660 45220
rect 30828 45052 30884 45108
rect 30492 42924 30548 42980
rect 30156 41244 30212 41300
rect 28476 40460 28532 40516
rect 27356 39564 27412 39620
rect 28364 40236 28420 40292
rect 27020 39004 27076 39060
rect 26684 37996 26740 38052
rect 26572 36988 26628 37044
rect 26572 36258 26628 36260
rect 26572 36206 26574 36258
rect 26574 36206 26626 36258
rect 26626 36206 26628 36258
rect 26572 36204 26628 36206
rect 27356 38220 27412 38276
rect 27356 37884 27412 37940
rect 26908 37212 26964 37268
rect 27244 37378 27300 37380
rect 27244 37326 27246 37378
rect 27246 37326 27298 37378
rect 27298 37326 27300 37378
rect 27244 37324 27300 37326
rect 26684 34748 26740 34804
rect 26908 35084 26964 35140
rect 26572 34018 26628 34020
rect 26572 33966 26574 34018
rect 26574 33966 26626 34018
rect 26626 33966 26628 34018
rect 26572 33964 26628 33966
rect 26236 32562 26292 32564
rect 26236 32510 26238 32562
rect 26238 32510 26290 32562
rect 26290 32510 26292 32562
rect 26236 32508 26292 32510
rect 26124 30156 26180 30212
rect 25676 29650 25732 29652
rect 25676 29598 25678 29650
rect 25678 29598 25730 29650
rect 25730 29598 25732 29650
rect 25676 29596 25732 29598
rect 29932 41020 29988 41076
rect 29708 40236 29764 40292
rect 27580 39058 27636 39060
rect 27580 39006 27582 39058
rect 27582 39006 27634 39058
rect 27634 39006 27636 39058
rect 27580 39004 27636 39006
rect 27804 38332 27860 38388
rect 28812 38332 28868 38388
rect 28812 37266 28868 37268
rect 28812 37214 28814 37266
rect 28814 37214 28866 37266
rect 28866 37214 28868 37266
rect 28812 37212 28868 37214
rect 29148 36988 29204 37044
rect 29708 36258 29764 36260
rect 29708 36206 29710 36258
rect 29710 36206 29762 36258
rect 29762 36206 29764 36258
rect 29708 36204 29764 36206
rect 29708 35810 29764 35812
rect 29708 35758 29710 35810
rect 29710 35758 29762 35810
rect 29762 35758 29764 35810
rect 29708 35756 29764 35758
rect 30044 40626 30100 40628
rect 30044 40574 30046 40626
rect 30046 40574 30098 40626
rect 30098 40574 30100 40626
rect 30044 40572 30100 40574
rect 30492 40460 30548 40516
rect 30044 36204 30100 36260
rect 30156 39004 30212 39060
rect 31164 45164 31220 45220
rect 31500 45388 31556 45444
rect 31388 44882 31444 44884
rect 31388 44830 31390 44882
rect 31390 44830 31442 44882
rect 31442 44830 31444 44882
rect 31388 44828 31444 44830
rect 31052 44322 31108 44324
rect 31052 44270 31054 44322
rect 31054 44270 31106 44322
rect 31106 44270 31108 44322
rect 31052 44268 31108 44270
rect 31724 46956 31780 47012
rect 38444 54684 38500 54740
rect 35980 54348 36036 54404
rect 35868 49922 35924 49924
rect 35868 49870 35870 49922
rect 35870 49870 35922 49922
rect 35922 49870 35924 49922
rect 35868 49868 35924 49870
rect 41132 56140 41188 56196
rect 42140 56194 42196 56196
rect 42140 56142 42142 56194
rect 42142 56142 42194 56194
rect 42194 56142 42196 56194
rect 42140 56140 42196 56142
rect 44940 56140 44996 56196
rect 40348 55356 40404 55412
rect 41244 55356 41300 55412
rect 42588 56028 42644 56084
rect 40348 54572 40404 54628
rect 39228 53842 39284 53844
rect 39228 53790 39230 53842
rect 39230 53790 39282 53842
rect 39282 53790 39284 53842
rect 39228 53788 39284 53790
rect 42364 53842 42420 53844
rect 42364 53790 42366 53842
rect 42366 53790 42418 53842
rect 42418 53790 42420 53842
rect 42364 53788 42420 53790
rect 39116 53506 39172 53508
rect 39116 53454 39118 53506
rect 39118 53454 39170 53506
rect 39170 53454 39172 53506
rect 39116 53452 39172 53454
rect 39564 53452 39620 53508
rect 37548 51212 37604 51268
rect 36764 50428 36820 50484
rect 35868 49138 35924 49140
rect 35868 49086 35870 49138
rect 35870 49086 35922 49138
rect 35922 49086 35924 49138
rect 35868 49084 35924 49086
rect 33852 48636 33908 48692
rect 32956 46562 33012 46564
rect 32956 46510 32958 46562
rect 32958 46510 33010 46562
rect 33010 46510 33012 46562
rect 32956 46508 33012 46510
rect 31724 45388 31780 45444
rect 31612 44380 31668 44436
rect 31948 45164 32004 45220
rect 32172 45218 32228 45220
rect 32172 45166 32174 45218
rect 32174 45166 32226 45218
rect 32226 45166 32228 45218
rect 32172 45164 32228 45166
rect 32620 45164 32676 45220
rect 32060 44716 32116 44772
rect 31276 43596 31332 43652
rect 31612 43650 31668 43652
rect 31612 43598 31614 43650
rect 31614 43598 31666 43650
rect 31666 43598 31668 43650
rect 31612 43596 31668 43598
rect 31500 43036 31556 43092
rect 31612 42140 31668 42196
rect 31388 42028 31444 42084
rect 31052 40572 31108 40628
rect 31164 40514 31220 40516
rect 31164 40462 31166 40514
rect 31166 40462 31218 40514
rect 31218 40462 31220 40514
rect 31164 40460 31220 40462
rect 30492 38220 30548 38276
rect 31276 39506 31332 39508
rect 31276 39454 31278 39506
rect 31278 39454 31330 39506
rect 31330 39454 31332 39506
rect 31276 39452 31332 39454
rect 30940 39058 30996 39060
rect 30940 39006 30942 39058
rect 30942 39006 30994 39058
rect 30994 39006 30996 39058
rect 30940 39004 30996 39006
rect 29932 35756 29988 35812
rect 29372 35196 29428 35252
rect 27916 34412 27972 34468
rect 27916 33964 27972 34020
rect 26796 32956 26852 33012
rect 26908 32732 26964 32788
rect 27804 33234 27860 33236
rect 27804 33182 27806 33234
rect 27806 33182 27858 33234
rect 27858 33182 27860 33234
rect 27804 33180 27860 33182
rect 27244 32844 27300 32900
rect 27692 33122 27748 33124
rect 27692 33070 27694 33122
rect 27694 33070 27746 33122
rect 27746 33070 27748 33122
rect 27692 33068 27748 33070
rect 27468 32956 27524 33012
rect 28476 34412 28532 34468
rect 28476 33740 28532 33796
rect 28028 33180 28084 33236
rect 27244 32620 27300 32676
rect 27580 32620 27636 32676
rect 25676 28924 25732 28980
rect 25228 26908 25284 26964
rect 23548 24892 23604 24948
rect 22428 24780 22484 24836
rect 22428 24610 22484 24612
rect 22428 24558 22430 24610
rect 22430 24558 22482 24610
rect 22482 24558 22484 24610
rect 22428 24556 22484 24558
rect 22764 24556 22820 24612
rect 22316 23772 22372 23828
rect 23212 23826 23268 23828
rect 23212 23774 23214 23826
rect 23214 23774 23266 23826
rect 23266 23774 23268 23826
rect 23212 23772 23268 23774
rect 23100 23660 23156 23716
rect 22988 23548 23044 23604
rect 21980 22988 22036 23044
rect 23660 25116 23716 25172
rect 24108 25282 24164 25284
rect 24108 25230 24110 25282
rect 24110 25230 24162 25282
rect 24162 25230 24164 25282
rect 24108 25228 24164 25230
rect 24668 25116 24724 25172
rect 23996 24668 24052 24724
rect 24108 25004 24164 25060
rect 23660 24610 23716 24612
rect 23660 24558 23662 24610
rect 23662 24558 23714 24610
rect 23714 24558 23716 24610
rect 23660 24556 23716 24558
rect 23548 23548 23604 23604
rect 22764 22988 22820 23044
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 12348 4508 12404 4564
rect 16492 5292 16548 5348
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 11788 3612 11844 3668
rect 8876 3388 8932 3444
rect 9996 3442 10052 3444
rect 9996 3390 9998 3442
rect 9998 3390 10050 3442
rect 10050 3390 10052 3442
rect 9996 3388 10052 3390
rect 16828 3666 16884 3668
rect 16828 3614 16830 3666
rect 16830 3614 16882 3666
rect 16882 3614 16884 3666
rect 16828 3612 16884 3614
rect 17724 3612 17780 3668
rect 20748 3442 20804 3444
rect 20748 3390 20750 3442
rect 20750 3390 20802 3442
rect 20802 3390 20804 3442
rect 20748 3388 20804 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21420 3442 21476 3444
rect 21420 3390 21422 3442
rect 21422 3390 21474 3442
rect 21474 3390 21476 3442
rect 21420 3388 21476 3390
rect 21756 3330 21812 3332
rect 21756 3278 21758 3330
rect 21758 3278 21810 3330
rect 21810 3278 21812 3330
rect 21756 3276 21812 3278
rect 24332 24892 24388 24948
rect 24220 24722 24276 24724
rect 24220 24670 24222 24722
rect 24222 24670 24274 24722
rect 24274 24670 24276 24722
rect 24220 24668 24276 24670
rect 24220 23996 24276 24052
rect 24668 24946 24724 24948
rect 24668 24894 24670 24946
rect 24670 24894 24722 24946
rect 24722 24894 24724 24946
rect 24668 24892 24724 24894
rect 26460 28924 26516 28980
rect 26908 30044 26964 30100
rect 26460 28754 26516 28756
rect 26460 28702 26462 28754
rect 26462 28702 26514 28754
rect 26514 28702 26516 28754
rect 26460 28700 26516 28702
rect 26908 28700 26964 28756
rect 25676 27132 25732 27188
rect 24444 24556 24500 24612
rect 24332 24108 24388 24164
rect 26012 27244 26068 27300
rect 26460 26962 26516 26964
rect 26460 26910 26462 26962
rect 26462 26910 26514 26962
rect 26514 26910 26516 26962
rect 26460 26908 26516 26910
rect 27244 32060 27300 32116
rect 27132 27468 27188 27524
rect 27020 27244 27076 27300
rect 27468 28700 27524 28756
rect 27692 27074 27748 27076
rect 27692 27022 27694 27074
rect 27694 27022 27746 27074
rect 27746 27022 27748 27074
rect 27692 27020 27748 27022
rect 28252 33234 28308 33236
rect 28252 33182 28254 33234
rect 28254 33182 28306 33234
rect 28306 33182 28308 33234
rect 28252 33180 28308 33182
rect 28924 33180 28980 33236
rect 28588 32844 28644 32900
rect 28924 32508 28980 32564
rect 30380 37938 30436 37940
rect 30380 37886 30382 37938
rect 30382 37886 30434 37938
rect 30434 37886 30436 37938
rect 30380 37884 30436 37886
rect 30940 37378 30996 37380
rect 30940 37326 30942 37378
rect 30942 37326 30994 37378
rect 30994 37326 30996 37378
rect 30940 37324 30996 37326
rect 31724 40908 31780 40964
rect 32060 43650 32116 43652
rect 32060 43598 32062 43650
rect 32062 43598 32114 43650
rect 32114 43598 32116 43650
rect 32060 43596 32116 43598
rect 32396 43260 32452 43316
rect 31836 40460 31892 40516
rect 32060 40626 32116 40628
rect 32060 40574 32062 40626
rect 32062 40574 32114 40626
rect 32114 40574 32116 40626
rect 32060 40572 32116 40574
rect 31836 40290 31892 40292
rect 31836 40238 31838 40290
rect 31838 40238 31890 40290
rect 31890 40238 31892 40290
rect 31836 40236 31892 40238
rect 31948 38892 32004 38948
rect 31500 38050 31556 38052
rect 31500 37998 31502 38050
rect 31502 37998 31554 38050
rect 31554 37998 31556 38050
rect 31500 37996 31556 37998
rect 31948 37884 32004 37940
rect 31276 37324 31332 37380
rect 30604 36482 30660 36484
rect 30604 36430 30606 36482
rect 30606 36430 30658 36482
rect 30658 36430 30660 36482
rect 30604 36428 30660 36430
rect 30380 36258 30436 36260
rect 30380 36206 30382 36258
rect 30382 36206 30434 36258
rect 30434 36206 30436 36258
rect 30380 36204 30436 36206
rect 30716 35756 30772 35812
rect 31500 37378 31556 37380
rect 31500 37326 31502 37378
rect 31502 37326 31554 37378
rect 31554 37326 31556 37378
rect 31500 37324 31556 37326
rect 32284 39506 32340 39508
rect 32284 39454 32286 39506
rect 32286 39454 32338 39506
rect 32338 39454 32340 39506
rect 32284 39452 32340 39454
rect 32060 37436 32116 37492
rect 32620 43372 32676 43428
rect 33740 46562 33796 46564
rect 33740 46510 33742 46562
rect 33742 46510 33794 46562
rect 33794 46510 33796 46562
rect 33740 46508 33796 46510
rect 33628 45276 33684 45332
rect 33516 44434 33572 44436
rect 33516 44382 33518 44434
rect 33518 44382 33570 44434
rect 33570 44382 33572 44434
rect 33516 44380 33572 44382
rect 33628 44268 33684 44324
rect 33068 43596 33124 43652
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34076 45778 34132 45780
rect 34076 45726 34078 45778
rect 34078 45726 34130 45778
rect 34130 45726 34132 45778
rect 34076 45724 34132 45726
rect 33964 44156 34020 44212
rect 34076 44268 34132 44324
rect 32956 43260 33012 43316
rect 33740 42028 33796 42084
rect 32620 41692 32676 41748
rect 34188 43596 34244 43652
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35644 45836 35700 45892
rect 34524 45778 34580 45780
rect 34524 45726 34526 45778
rect 34526 45726 34578 45778
rect 34578 45726 34580 45778
rect 34524 45724 34580 45726
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34300 43484 34356 43540
rect 34188 43372 34244 43428
rect 35084 43314 35140 43316
rect 35084 43262 35086 43314
rect 35086 43262 35138 43314
rect 35138 43262 35140 43314
rect 35084 43260 35140 43262
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35420 41692 35476 41748
rect 35532 41804 35588 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35980 45500 36036 45556
rect 36428 48802 36484 48804
rect 36428 48750 36430 48802
rect 36430 48750 36482 48802
rect 36482 48750 36484 48802
rect 36428 48748 36484 48750
rect 36988 48748 37044 48804
rect 36652 45836 36708 45892
rect 36764 48300 36820 48356
rect 36652 44940 36708 44996
rect 35644 41468 35700 41524
rect 37436 48802 37492 48804
rect 37436 48750 37438 48802
rect 37438 48750 37490 48802
rect 37490 48750 37492 48802
rect 37436 48748 37492 48750
rect 37100 45836 37156 45892
rect 38556 51266 38612 51268
rect 38556 51214 38558 51266
rect 38558 51214 38610 51266
rect 38610 51214 38612 51266
rect 38556 51212 38612 51214
rect 39452 50988 39508 51044
rect 37772 49756 37828 49812
rect 36988 45724 37044 45780
rect 37324 45218 37380 45220
rect 37324 45166 37326 45218
rect 37326 45166 37378 45218
rect 37378 45166 37380 45218
rect 37324 45164 37380 45166
rect 36988 44940 37044 44996
rect 35532 41356 35588 41412
rect 35308 41244 35364 41300
rect 33404 40962 33460 40964
rect 33404 40910 33406 40962
rect 33406 40910 33458 40962
rect 33458 40910 33460 40962
rect 33404 40908 33460 40910
rect 32620 40626 32676 40628
rect 32620 40574 32622 40626
rect 32622 40574 32674 40626
rect 32674 40574 32676 40626
rect 32620 40572 32676 40574
rect 32508 38108 32564 38164
rect 33068 40236 33124 40292
rect 32844 38050 32900 38052
rect 32844 37998 32846 38050
rect 32846 37998 32898 38050
rect 32898 37998 32900 38050
rect 32844 37996 32900 37998
rect 31948 37100 32004 37156
rect 32284 36764 32340 36820
rect 31388 36428 31444 36484
rect 32172 36482 32228 36484
rect 32172 36430 32174 36482
rect 32174 36430 32226 36482
rect 32226 36430 32228 36482
rect 32172 36428 32228 36430
rect 32620 37490 32676 37492
rect 32620 37438 32622 37490
rect 32622 37438 32674 37490
rect 32674 37438 32676 37490
rect 32620 37436 32676 37438
rect 32732 36764 32788 36820
rect 32396 35698 32452 35700
rect 32396 35646 32398 35698
rect 32398 35646 32450 35698
rect 32450 35646 32452 35698
rect 32396 35644 32452 35646
rect 32844 35532 32900 35588
rect 31500 35420 31556 35476
rect 30156 35196 30212 35252
rect 29596 35138 29652 35140
rect 29596 35086 29598 35138
rect 29598 35086 29650 35138
rect 29650 35086 29652 35138
rect 29596 35084 29652 35086
rect 29484 34524 29540 34580
rect 29708 34076 29764 34132
rect 33180 40012 33236 40068
rect 35084 41020 35140 41076
rect 34636 40908 34692 40964
rect 33852 40348 33908 40404
rect 34300 40236 34356 40292
rect 34076 40124 34132 40180
rect 33180 39228 33236 39284
rect 33180 37436 33236 37492
rect 33180 36988 33236 37044
rect 33516 36652 33572 36708
rect 33516 36482 33572 36484
rect 33516 36430 33518 36482
rect 33518 36430 33570 36482
rect 33570 36430 33572 36482
rect 33516 36428 33572 36430
rect 33740 39228 33796 39284
rect 33964 38050 34020 38052
rect 33964 37998 33966 38050
rect 33966 37998 34018 38050
rect 34018 37998 34020 38050
rect 33964 37996 34020 37998
rect 33964 37212 34020 37268
rect 34524 39900 34580 39956
rect 34860 40626 34916 40628
rect 34860 40574 34862 40626
rect 34862 40574 34914 40626
rect 34914 40574 34916 40626
rect 34860 40572 34916 40574
rect 35084 40460 35140 40516
rect 34972 40348 35028 40404
rect 34748 40178 34804 40180
rect 34748 40126 34750 40178
rect 34750 40126 34802 40178
rect 34802 40126 34804 40178
rect 34748 40124 34804 40126
rect 34636 39788 34692 39844
rect 34524 39340 34580 39396
rect 36876 43650 36932 43652
rect 36876 43598 36878 43650
rect 36878 43598 36930 43650
rect 36930 43598 36932 43650
rect 36876 43596 36932 43598
rect 36652 43538 36708 43540
rect 36652 43486 36654 43538
rect 36654 43486 36706 43538
rect 36706 43486 36708 43538
rect 36652 43484 36708 43486
rect 35980 43426 36036 43428
rect 35980 43374 35982 43426
rect 35982 43374 36034 43426
rect 36034 43374 36036 43426
rect 35980 43372 36036 43374
rect 36204 42530 36260 42532
rect 36204 42478 36206 42530
rect 36206 42478 36258 42530
rect 36258 42478 36260 42530
rect 36204 42476 36260 42478
rect 36652 42476 36708 42532
rect 37100 43426 37156 43428
rect 37100 43374 37102 43426
rect 37102 43374 37154 43426
rect 37154 43374 37156 43426
rect 37100 43372 37156 43374
rect 36428 41298 36484 41300
rect 36428 41246 36430 41298
rect 36430 41246 36482 41298
rect 36482 41246 36484 41298
rect 36428 41244 36484 41246
rect 35980 41074 36036 41076
rect 35980 41022 35982 41074
rect 35982 41022 36034 41074
rect 36034 41022 36036 41074
rect 35980 41020 36036 41022
rect 35980 40572 36036 40628
rect 36204 40460 36260 40516
rect 35980 40402 36036 40404
rect 35980 40350 35982 40402
rect 35982 40350 36034 40402
rect 36034 40350 36036 40402
rect 35980 40348 36036 40350
rect 36540 40348 36596 40404
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35644 40012 35700 40068
rect 35084 39618 35140 39620
rect 35084 39566 35086 39618
rect 35086 39566 35138 39618
rect 35138 39566 35140 39618
rect 35084 39564 35140 39566
rect 36428 39676 36484 39732
rect 35084 39340 35140 39396
rect 35756 39394 35812 39396
rect 35756 39342 35758 39394
rect 35758 39342 35810 39394
rect 35810 39342 35812 39394
rect 35756 39340 35812 39342
rect 35644 39228 35700 39284
rect 35756 39116 35812 39172
rect 33628 35980 33684 36036
rect 33180 35756 33236 35812
rect 33628 35810 33684 35812
rect 33628 35758 33630 35810
rect 33630 35758 33682 35810
rect 33682 35758 33684 35810
rect 33628 35756 33684 35758
rect 34076 36706 34132 36708
rect 34076 36654 34078 36706
rect 34078 36654 34130 36706
rect 34130 36654 34132 36706
rect 34076 36652 34132 36654
rect 36204 39116 36260 39172
rect 35868 38556 35924 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34412 38162 34468 38164
rect 34412 38110 34414 38162
rect 34414 38110 34466 38162
rect 34466 38110 34468 38162
rect 34412 38108 34468 38110
rect 35084 38162 35140 38164
rect 35084 38110 35086 38162
rect 35086 38110 35138 38162
rect 35138 38110 35140 38162
rect 35084 38108 35140 38110
rect 35308 38050 35364 38052
rect 35308 37998 35310 38050
rect 35310 37998 35362 38050
rect 35362 37998 35364 38050
rect 35308 37996 35364 37998
rect 35084 37100 35140 37156
rect 34972 36652 35028 36708
rect 34076 36482 34132 36484
rect 34076 36430 34078 36482
rect 34078 36430 34130 36482
rect 34130 36430 34132 36482
rect 34076 36428 34132 36430
rect 34412 36594 34468 36596
rect 34412 36542 34414 36594
rect 34414 36542 34466 36594
rect 34466 36542 34468 36594
rect 34412 36540 34468 36542
rect 33740 35532 33796 35588
rect 33852 34076 33908 34132
rect 29708 33404 29764 33460
rect 29596 33234 29652 33236
rect 29596 33182 29598 33234
rect 29598 33182 29650 33234
rect 29650 33182 29652 33234
rect 29596 33180 29652 33182
rect 30268 33458 30324 33460
rect 30268 33406 30270 33458
rect 30270 33406 30322 33458
rect 30322 33406 30324 33458
rect 30268 33404 30324 33406
rect 29372 32284 29428 32340
rect 29484 32956 29540 33012
rect 28140 31836 28196 31892
rect 30492 31890 30548 31892
rect 30492 31838 30494 31890
rect 30494 31838 30546 31890
rect 30546 31838 30548 31890
rect 30492 31836 30548 31838
rect 29932 31724 29988 31780
rect 30604 31388 30660 31444
rect 30828 31164 30884 31220
rect 31724 31388 31780 31444
rect 31276 31164 31332 31220
rect 28028 30044 28084 30100
rect 28700 30882 28756 30884
rect 28700 30830 28702 30882
rect 28702 30830 28754 30882
rect 28754 30830 28756 30882
rect 28700 30828 28756 30830
rect 28028 28812 28084 28868
rect 27916 28754 27972 28756
rect 27916 28702 27918 28754
rect 27918 28702 27970 28754
rect 27970 28702 27972 28754
rect 27916 28700 27972 28702
rect 28028 28588 28084 28644
rect 27132 26796 27188 26852
rect 26908 25004 26964 25060
rect 27916 27692 27972 27748
rect 27916 27132 27972 27188
rect 27244 26514 27300 26516
rect 27244 26462 27246 26514
rect 27246 26462 27298 26514
rect 27298 26462 27300 26514
rect 27244 26460 27300 26462
rect 27804 26514 27860 26516
rect 27804 26462 27806 26514
rect 27806 26462 27858 26514
rect 27858 26462 27860 26514
rect 27804 26460 27860 26462
rect 27132 25004 27188 25060
rect 27468 24946 27524 24948
rect 27468 24894 27470 24946
rect 27470 24894 27522 24946
rect 27522 24894 27524 24946
rect 27468 24892 27524 24894
rect 27916 24780 27972 24836
rect 26348 24108 26404 24164
rect 24220 23660 24276 23716
rect 28924 29260 28980 29316
rect 28476 29148 28532 29204
rect 28476 28754 28532 28756
rect 28476 28702 28478 28754
rect 28478 28702 28530 28754
rect 28530 28702 28532 28754
rect 28476 28700 28532 28702
rect 28252 27020 28308 27076
rect 28812 28700 28868 28756
rect 28588 28476 28644 28532
rect 28700 28082 28756 28084
rect 28700 28030 28702 28082
rect 28702 28030 28754 28082
rect 28754 28030 28756 28082
rect 28700 28028 28756 28030
rect 28700 27634 28756 27636
rect 28700 27582 28702 27634
rect 28702 27582 28754 27634
rect 28754 27582 28756 27634
rect 28700 27580 28756 27582
rect 28588 27244 28644 27300
rect 28700 27020 28756 27076
rect 28364 25004 28420 25060
rect 29260 28476 29316 28532
rect 31164 28476 31220 28532
rect 31612 29986 31668 29988
rect 31612 29934 31614 29986
rect 31614 29934 31666 29986
rect 31666 29934 31668 29986
rect 31612 29932 31668 29934
rect 29260 28082 29316 28084
rect 29260 28030 29262 28082
rect 29262 28030 29314 28082
rect 29314 28030 29316 28082
rect 29260 28028 29316 28030
rect 29484 27244 29540 27300
rect 31276 27186 31332 27188
rect 31276 27134 31278 27186
rect 31278 27134 31330 27186
rect 31330 27134 31332 27186
rect 31276 27132 31332 27134
rect 31612 27132 31668 27188
rect 31724 27074 31780 27076
rect 31724 27022 31726 27074
rect 31726 27022 31778 27074
rect 31778 27022 31780 27074
rect 31724 27020 31780 27022
rect 28924 25004 28980 25060
rect 28588 24946 28644 24948
rect 28588 24894 28590 24946
rect 28590 24894 28642 24946
rect 28642 24894 28644 24946
rect 28588 24892 28644 24894
rect 28812 24834 28868 24836
rect 28812 24782 28814 24834
rect 28814 24782 28866 24834
rect 28866 24782 28868 24834
rect 28812 24780 28868 24782
rect 28812 11116 28868 11172
rect 32508 32956 32564 33012
rect 33068 32956 33124 33012
rect 32060 32396 32116 32452
rect 34076 33516 34132 33572
rect 34188 35644 34244 35700
rect 33964 32786 34020 32788
rect 33964 32734 33966 32786
rect 33966 32734 34018 32786
rect 34018 32734 34020 32786
rect 33964 32732 34020 32734
rect 34860 36594 34916 36596
rect 34860 36542 34862 36594
rect 34862 36542 34914 36594
rect 34914 36542 34916 36594
rect 34860 36540 34916 36542
rect 34636 36428 34692 36484
rect 34412 35698 34468 35700
rect 34412 35646 34414 35698
rect 34414 35646 34466 35698
rect 34466 35646 34468 35698
rect 34412 35644 34468 35646
rect 34860 35980 34916 36036
rect 34972 35756 35028 35812
rect 36092 38668 36148 38724
rect 35868 36988 35924 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 36540 35588 36596
rect 35196 35306 35252 35308
rect 34972 35196 35028 35252
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35644 35810 35700 35812
rect 35644 35758 35646 35810
rect 35646 35758 35698 35810
rect 35698 35758 35700 35810
rect 35644 35756 35700 35758
rect 35980 36428 36036 36484
rect 35980 35980 36036 36036
rect 35756 35532 35812 35588
rect 34636 34130 34692 34132
rect 34636 34078 34638 34130
rect 34638 34078 34690 34130
rect 34690 34078 34692 34130
rect 34636 34076 34692 34078
rect 35084 34636 35140 34692
rect 34860 33516 34916 33572
rect 34972 34300 35028 34356
rect 34524 32786 34580 32788
rect 34524 32734 34526 32786
rect 34526 32734 34578 32786
rect 34578 32734 34580 32786
rect 34524 32732 34580 32734
rect 33628 30156 33684 30212
rect 32172 29986 32228 29988
rect 32172 29934 32174 29986
rect 32174 29934 32226 29986
rect 32226 29934 32228 29986
rect 32172 29932 32228 29934
rect 32172 29314 32228 29316
rect 32172 29262 32174 29314
rect 32174 29262 32226 29314
rect 32226 29262 32228 29314
rect 32172 29260 32228 29262
rect 32732 29314 32788 29316
rect 32732 29262 32734 29314
rect 32734 29262 32786 29314
rect 32786 29262 32788 29314
rect 32732 29260 32788 29262
rect 32620 28700 32676 28756
rect 33292 28812 33348 28868
rect 33628 28812 33684 28868
rect 33740 28700 33796 28756
rect 32844 28588 32900 28644
rect 32396 28476 32452 28532
rect 32732 27692 32788 27748
rect 32732 27074 32788 27076
rect 32732 27022 32734 27074
rect 32734 27022 32786 27074
rect 32786 27022 32788 27074
rect 32732 27020 32788 27022
rect 33292 27132 33348 27188
rect 33964 27244 34020 27300
rect 34076 28252 34132 28308
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35420 33346 35476 33348
rect 35420 33294 35422 33346
rect 35422 33294 35474 33346
rect 35474 33294 35476 33346
rect 35420 33292 35476 33294
rect 35644 33292 35700 33348
rect 35196 32732 35252 32788
rect 35532 33068 35588 33124
rect 35868 35308 35924 35364
rect 36652 40290 36708 40292
rect 36652 40238 36654 40290
rect 36654 40238 36706 40290
rect 36706 40238 36708 40290
rect 36652 40236 36708 40238
rect 36540 39340 36596 39396
rect 36316 38892 36372 38948
rect 36204 37490 36260 37492
rect 36204 37438 36206 37490
rect 36206 37438 36258 37490
rect 36258 37438 36260 37490
rect 36204 37436 36260 37438
rect 36316 35308 36372 35364
rect 35868 34300 35924 34356
rect 36316 35084 36372 35140
rect 35196 32396 35252 32452
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35868 32450 35924 32452
rect 35868 32398 35870 32450
rect 35870 32398 35922 32450
rect 35922 32398 35924 32450
rect 35868 32396 35924 32398
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34524 29260 34580 29316
rect 35756 29260 35812 29316
rect 35196 29034 35252 29036
rect 34636 28924 34692 28980
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35756 28924 35812 28980
rect 34636 28754 34692 28756
rect 34636 28702 34638 28754
rect 34638 28702 34690 28754
rect 34690 28702 34692 28754
rect 34636 28700 34692 28702
rect 35308 28812 35364 28868
rect 35308 28588 35364 28644
rect 35532 28700 35588 28756
rect 36092 34690 36148 34692
rect 36092 34638 36094 34690
rect 36094 34638 36146 34690
rect 36146 34638 36148 34690
rect 36092 34636 36148 34638
rect 36092 34354 36148 34356
rect 36092 34302 36094 34354
rect 36094 34302 36146 34354
rect 36146 34302 36148 34354
rect 36092 34300 36148 34302
rect 36092 33068 36148 33124
rect 36652 38556 36708 38612
rect 36652 37436 36708 37492
rect 36540 36540 36596 36596
rect 36652 35532 36708 35588
rect 36652 35308 36708 35364
rect 36428 33404 36484 33460
rect 36204 31388 36260 31444
rect 36876 41468 36932 41524
rect 36876 34860 36932 34916
rect 36764 33964 36820 34020
rect 36652 33180 36708 33236
rect 35420 28418 35476 28420
rect 35420 28366 35422 28418
rect 35422 28366 35474 28418
rect 35474 28366 35476 28418
rect 35420 28364 35476 28366
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 39452 50482 39508 50484
rect 39452 50430 39454 50482
rect 39454 50430 39506 50482
rect 39506 50430 39508 50482
rect 39452 50428 39508 50430
rect 39004 48636 39060 48692
rect 37996 48076 38052 48132
rect 38556 48130 38612 48132
rect 38556 48078 38558 48130
rect 38558 48078 38610 48130
rect 38610 48078 38612 48130
rect 38556 48076 38612 48078
rect 38332 47068 38388 47124
rect 37884 45666 37940 45668
rect 37884 45614 37886 45666
rect 37886 45614 37938 45666
rect 37938 45614 37940 45666
rect 37884 45612 37940 45614
rect 37996 45890 38052 45892
rect 37996 45838 37998 45890
rect 37998 45838 38050 45890
rect 38050 45838 38052 45890
rect 37996 45836 38052 45838
rect 37772 44994 37828 44996
rect 37772 44942 37774 44994
rect 37774 44942 37826 44994
rect 37826 44942 37828 44994
rect 37772 44940 37828 44942
rect 37660 43484 37716 43540
rect 39004 45666 39060 45668
rect 39004 45614 39006 45666
rect 39006 45614 39058 45666
rect 39058 45614 39060 45666
rect 39004 45612 39060 45614
rect 38556 45276 38612 45332
rect 38220 45218 38276 45220
rect 38220 45166 38222 45218
rect 38222 45166 38274 45218
rect 38274 45166 38276 45218
rect 38220 45164 38276 45166
rect 40012 53506 40068 53508
rect 40012 53454 40014 53506
rect 40014 53454 40066 53506
rect 40066 53454 40068 53506
rect 40012 53452 40068 53454
rect 40684 53506 40740 53508
rect 40684 53454 40686 53506
rect 40686 53454 40738 53506
rect 40738 53454 40740 53506
rect 40684 53452 40740 53454
rect 40796 53340 40852 53396
rect 39900 52108 39956 52164
rect 40236 51436 40292 51492
rect 39900 51212 39956 51268
rect 40684 51324 40740 51380
rect 40796 52108 40852 52164
rect 41692 53506 41748 53508
rect 41692 53454 41694 53506
rect 41694 53454 41746 53506
rect 41746 53454 41748 53506
rect 41692 53452 41748 53454
rect 41468 53340 41524 53396
rect 41244 51548 41300 51604
rect 42140 53564 42196 53620
rect 41468 51436 41524 51492
rect 42476 51324 42532 51380
rect 40236 50988 40292 51044
rect 40012 50764 40068 50820
rect 40460 50818 40516 50820
rect 40460 50766 40462 50818
rect 40462 50766 40514 50818
rect 40514 50766 40516 50818
rect 40460 50764 40516 50766
rect 40124 47068 40180 47124
rect 40236 50482 40292 50484
rect 40236 50430 40238 50482
rect 40238 50430 40290 50482
rect 40290 50430 40292 50482
rect 40236 50428 40292 50430
rect 40908 50482 40964 50484
rect 40908 50430 40910 50482
rect 40910 50430 40962 50482
rect 40962 50430 40964 50482
rect 40908 50428 40964 50430
rect 39900 45330 39956 45332
rect 39900 45278 39902 45330
rect 39902 45278 39954 45330
rect 39954 45278 39956 45330
rect 39900 45276 39956 45278
rect 40012 44994 40068 44996
rect 40012 44942 40014 44994
rect 40014 44942 40066 44994
rect 40066 44942 40068 44994
rect 40012 44940 40068 44942
rect 42140 51100 42196 51156
rect 42476 48076 42532 48132
rect 41580 46396 41636 46452
rect 41804 46620 41860 46676
rect 41020 45724 41076 45780
rect 40796 45388 40852 45444
rect 37996 43372 38052 43428
rect 37324 43314 37380 43316
rect 37324 43262 37326 43314
rect 37326 43262 37378 43314
rect 37378 43262 37380 43314
rect 37324 43260 37380 43262
rect 37548 41580 37604 41636
rect 37660 42812 37716 42868
rect 37660 41244 37716 41300
rect 37884 41916 37940 41972
rect 37548 40962 37604 40964
rect 37548 40910 37550 40962
rect 37550 40910 37602 40962
rect 37602 40910 37604 40962
rect 37548 40908 37604 40910
rect 39676 41692 39732 41748
rect 39228 41020 39284 41076
rect 37884 40796 37940 40852
rect 38556 40908 38612 40964
rect 38556 40572 38612 40628
rect 38780 40796 38836 40852
rect 38780 40348 38836 40404
rect 37548 40012 37604 40068
rect 38556 39788 38612 39844
rect 38332 39730 38388 39732
rect 38332 39678 38334 39730
rect 38334 39678 38386 39730
rect 38386 39678 38388 39730
rect 38332 39676 38388 39678
rect 38108 39618 38164 39620
rect 38108 39566 38110 39618
rect 38110 39566 38162 39618
rect 38162 39566 38164 39618
rect 38108 39564 38164 39566
rect 38780 39506 38836 39508
rect 38780 39454 38782 39506
rect 38782 39454 38834 39506
rect 38834 39454 38836 39506
rect 38780 39452 38836 39454
rect 39228 39506 39284 39508
rect 39228 39454 39230 39506
rect 39230 39454 39282 39506
rect 39282 39454 39284 39506
rect 39228 39452 39284 39454
rect 39116 38946 39172 38948
rect 39116 38894 39118 38946
rect 39118 38894 39170 38946
rect 39170 38894 39172 38946
rect 39116 38892 39172 38894
rect 38556 38668 38612 38724
rect 37212 36540 37268 36596
rect 38444 37884 38500 37940
rect 37100 36316 37156 36372
rect 37436 36316 37492 36372
rect 36988 34412 37044 34468
rect 37100 35756 37156 35812
rect 36988 34018 37044 34020
rect 36988 33966 36990 34018
rect 36990 33966 37042 34018
rect 37042 33966 37044 34018
rect 36988 33964 37044 33966
rect 38220 35810 38276 35812
rect 38220 35758 38222 35810
rect 38222 35758 38274 35810
rect 38274 35758 38276 35810
rect 38220 35756 38276 35758
rect 38108 35420 38164 35476
rect 37100 32844 37156 32900
rect 37324 33180 37380 33236
rect 37212 32786 37268 32788
rect 37212 32734 37214 32786
rect 37214 32734 37266 32786
rect 37266 32734 37268 32786
rect 37212 32732 37268 32734
rect 36988 32396 37044 32452
rect 36876 31778 36932 31780
rect 36876 31726 36878 31778
rect 36878 31726 36930 31778
rect 36930 31726 36932 31778
rect 36876 31724 36932 31726
rect 36988 30940 37044 30996
rect 37436 30156 37492 30212
rect 36764 28924 36820 28980
rect 37884 32732 37940 32788
rect 38332 33570 38388 33572
rect 38332 33518 38334 33570
rect 38334 33518 38386 33570
rect 38386 33518 38388 33570
rect 38332 33516 38388 33518
rect 38220 32956 38276 33012
rect 39116 37938 39172 37940
rect 39116 37886 39118 37938
rect 39118 37886 39170 37938
rect 39170 37886 39172 37938
rect 39116 37884 39172 37886
rect 38668 35586 38724 35588
rect 38668 35534 38670 35586
rect 38670 35534 38722 35586
rect 38722 35534 38724 35586
rect 38668 35532 38724 35534
rect 39116 35196 39172 35252
rect 39116 34412 39172 34468
rect 39900 41580 39956 41636
rect 40012 40908 40068 40964
rect 40236 40908 40292 40964
rect 40572 40908 40628 40964
rect 39900 39618 39956 39620
rect 39900 39566 39902 39618
rect 39902 39566 39954 39618
rect 39954 39566 39956 39618
rect 39900 39564 39956 39566
rect 40460 40684 40516 40740
rect 40236 40348 40292 40404
rect 40684 40796 40740 40852
rect 40796 40124 40852 40180
rect 40684 40012 40740 40068
rect 40572 39842 40628 39844
rect 40572 39790 40574 39842
rect 40574 39790 40626 39842
rect 40626 39790 40628 39842
rect 40572 39788 40628 39790
rect 40572 39564 40628 39620
rect 40684 39340 40740 39396
rect 40572 38946 40628 38948
rect 40572 38894 40574 38946
rect 40574 38894 40626 38946
rect 40626 38894 40628 38946
rect 40572 38892 40628 38894
rect 39452 37826 39508 37828
rect 39452 37774 39454 37826
rect 39454 37774 39506 37826
rect 39506 37774 39508 37826
rect 39452 37772 39508 37774
rect 39788 38050 39844 38052
rect 39788 37998 39790 38050
rect 39790 37998 39842 38050
rect 39842 37998 39844 38050
rect 39788 37996 39844 37998
rect 39788 36876 39844 36932
rect 39564 36258 39620 36260
rect 39564 36206 39566 36258
rect 39566 36206 39618 36258
rect 39618 36206 39620 36258
rect 39564 36204 39620 36206
rect 39676 36092 39732 36148
rect 39564 35810 39620 35812
rect 39564 35758 39566 35810
rect 39566 35758 39618 35810
rect 39618 35758 39620 35810
rect 39564 35756 39620 35758
rect 39788 35532 39844 35588
rect 40460 37212 40516 37268
rect 40124 36428 40180 36484
rect 40012 36370 40068 36372
rect 40012 36318 40014 36370
rect 40014 36318 40066 36370
rect 40066 36318 40068 36370
rect 40012 36316 40068 36318
rect 40012 35586 40068 35588
rect 40012 35534 40014 35586
rect 40014 35534 40066 35586
rect 40066 35534 40068 35586
rect 40012 35532 40068 35534
rect 40572 36652 40628 36708
rect 40908 38668 40964 38724
rect 40684 36258 40740 36260
rect 40684 36206 40686 36258
rect 40686 36206 40738 36258
rect 40738 36206 40740 36258
rect 40684 36204 40740 36206
rect 40236 35084 40292 35140
rect 39900 34188 39956 34244
rect 39228 33852 39284 33908
rect 38108 31778 38164 31780
rect 38108 31726 38110 31778
rect 38110 31726 38162 31778
rect 38162 31726 38164 31778
rect 38108 31724 38164 31726
rect 38444 32338 38500 32340
rect 38444 32286 38446 32338
rect 38446 32286 38498 32338
rect 38498 32286 38500 32338
rect 38444 32284 38500 32286
rect 38892 33180 38948 33236
rect 39004 32956 39060 33012
rect 39004 32060 39060 32116
rect 38668 31836 38724 31892
rect 39228 31890 39284 31892
rect 39228 31838 39230 31890
rect 39230 31838 39282 31890
rect 39282 31838 39284 31890
rect 39228 31836 39284 31838
rect 37772 31612 37828 31668
rect 37884 31500 37940 31556
rect 39452 31666 39508 31668
rect 39452 31614 39454 31666
rect 39454 31614 39506 31666
rect 39506 31614 39508 31666
rect 39452 31612 39508 31614
rect 39900 32620 39956 32676
rect 40124 32450 40180 32452
rect 40124 32398 40126 32450
rect 40126 32398 40178 32450
rect 40178 32398 40180 32450
rect 40124 32396 40180 32398
rect 39900 32060 39956 32116
rect 40012 31948 40068 32004
rect 39564 31500 39620 31556
rect 39900 31388 39956 31444
rect 40572 35196 40628 35252
rect 40348 31948 40404 32004
rect 40124 31388 40180 31444
rect 40348 31612 40404 31668
rect 40124 30882 40180 30884
rect 40124 30830 40126 30882
rect 40126 30830 40178 30882
rect 40178 30830 40180 30882
rect 40124 30828 40180 30830
rect 37996 30156 38052 30212
rect 37660 28700 37716 28756
rect 38108 29148 38164 29204
rect 39340 28812 39396 28868
rect 38108 28642 38164 28644
rect 38108 28590 38110 28642
rect 38110 28590 38162 28642
rect 38162 28590 38164 28642
rect 38108 28588 38164 28590
rect 36316 28252 36372 28308
rect 38556 28252 38612 28308
rect 39564 28642 39620 28644
rect 39564 28590 39566 28642
rect 39566 28590 39618 28642
rect 39618 28590 39620 28642
rect 39564 28588 39620 28590
rect 39900 28642 39956 28644
rect 39900 28590 39902 28642
rect 39902 28590 39954 28642
rect 39954 28590 39956 28642
rect 39900 28588 39956 28590
rect 39116 28252 39172 28308
rect 36092 27692 36148 27748
rect 35980 26908 36036 26964
rect 32508 23996 32564 24052
rect 28140 3276 28196 3332
rect 30156 3330 30212 3332
rect 30156 3278 30158 3330
rect 30158 3278 30210 3330
rect 30210 3278 30212 3330
rect 30156 3276 30212 3278
rect 39900 26348 39956 26404
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 40572 34076 40628 34132
rect 40908 33292 40964 33348
rect 40460 31500 40516 31556
rect 40684 32284 40740 32340
rect 40572 31388 40628 31444
rect 40460 28642 40516 28644
rect 40460 28590 40462 28642
rect 40462 28590 40514 28642
rect 40514 28590 40516 28642
rect 40460 28588 40516 28590
rect 40348 8092 40404 8148
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 31612 3276 31668 3332
rect 32396 3388 32452 3444
rect 34076 3442 34132 3444
rect 34076 3390 34078 3442
rect 34078 3390 34130 3442
rect 34130 3390 34132 3442
rect 34076 3388 34132 3390
rect 41244 44940 41300 44996
rect 41132 40684 41188 40740
rect 41132 38162 41188 38164
rect 41132 38110 41134 38162
rect 41134 38110 41186 38162
rect 41186 38110 41188 38162
rect 41132 38108 41188 38110
rect 41132 37100 41188 37156
rect 41132 36482 41188 36484
rect 41132 36430 41134 36482
rect 41134 36430 41186 36482
rect 41186 36430 41188 36482
rect 41132 36428 41188 36430
rect 41580 44994 41636 44996
rect 41580 44942 41582 44994
rect 41582 44942 41634 44994
rect 41634 44942 41636 44994
rect 41580 44940 41636 44942
rect 42364 46562 42420 46564
rect 42364 46510 42366 46562
rect 42366 46510 42418 46562
rect 42418 46510 42420 46562
rect 42364 46508 42420 46510
rect 41804 41916 41860 41972
rect 41916 45388 41972 45444
rect 41468 40402 41524 40404
rect 41468 40350 41470 40402
rect 41470 40350 41522 40402
rect 41522 40350 41524 40402
rect 41468 40348 41524 40350
rect 42812 53618 42868 53620
rect 42812 53566 42814 53618
rect 42814 53566 42866 53618
rect 42866 53566 42868 53618
rect 42812 53564 42868 53566
rect 42700 53058 42756 53060
rect 42700 53006 42702 53058
rect 42702 53006 42754 53058
rect 42754 53006 42756 53058
rect 42700 53004 42756 53006
rect 43372 53058 43428 53060
rect 43372 53006 43374 53058
rect 43374 53006 43426 53058
rect 43426 53006 43428 53058
rect 43372 53004 43428 53006
rect 43148 51100 43204 51156
rect 43036 50764 43092 50820
rect 43596 52834 43652 52836
rect 43596 52782 43598 52834
rect 43598 52782 43650 52834
rect 43650 52782 43652 52834
rect 43596 52780 43652 52782
rect 44044 52834 44100 52836
rect 44044 52782 44046 52834
rect 44046 52782 44098 52834
rect 44098 52782 44100 52834
rect 44044 52780 44100 52782
rect 43484 51378 43540 51380
rect 43484 51326 43486 51378
rect 43486 51326 43538 51378
rect 43538 51326 43540 51378
rect 43484 51324 43540 51326
rect 43596 50034 43652 50036
rect 43596 49982 43598 50034
rect 43598 49982 43650 50034
rect 43650 49982 43652 50034
rect 43596 49980 43652 49982
rect 43036 47964 43092 48020
rect 42924 46674 42980 46676
rect 42924 46622 42926 46674
rect 42926 46622 42978 46674
rect 42978 46622 42980 46674
rect 42924 46620 42980 46622
rect 43148 45388 43204 45444
rect 42812 41298 42868 41300
rect 42812 41246 42814 41298
rect 42814 41246 42866 41298
rect 42866 41246 42868 41298
rect 42812 41244 42868 41246
rect 41804 39788 41860 39844
rect 42028 40796 42084 40852
rect 42140 40684 42196 40740
rect 42700 40684 42756 40740
rect 42476 40236 42532 40292
rect 42812 39564 42868 39620
rect 41580 39394 41636 39396
rect 41580 39342 41582 39394
rect 41582 39342 41634 39394
rect 41634 39342 41636 39394
rect 41580 39340 41636 39342
rect 41916 38892 41972 38948
rect 41580 38722 41636 38724
rect 41580 38670 41582 38722
rect 41582 38670 41634 38722
rect 41634 38670 41636 38722
rect 41580 38668 41636 38670
rect 41692 38162 41748 38164
rect 41692 38110 41694 38162
rect 41694 38110 41746 38162
rect 41746 38110 41748 38162
rect 41692 38108 41748 38110
rect 41468 37266 41524 37268
rect 41468 37214 41470 37266
rect 41470 37214 41522 37266
rect 41522 37214 41524 37266
rect 41468 37212 41524 37214
rect 41692 36876 41748 36932
rect 41356 36706 41412 36708
rect 41356 36654 41358 36706
rect 41358 36654 41410 36706
rect 41410 36654 41412 36706
rect 41356 36652 41412 36654
rect 41580 36594 41636 36596
rect 41580 36542 41582 36594
rect 41582 36542 41634 36594
rect 41634 36542 41636 36594
rect 41580 36540 41636 36542
rect 42140 38050 42196 38052
rect 42140 37998 42142 38050
rect 42142 37998 42194 38050
rect 42194 37998 42196 38050
rect 42140 37996 42196 37998
rect 41916 36876 41972 36932
rect 42476 37436 42532 37492
rect 49532 56082 49588 56084
rect 49532 56030 49534 56082
rect 49534 56030 49586 56082
rect 49586 56030 49588 56082
rect 49532 56028 49588 56030
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 52780 56194 52836 56196
rect 52780 56142 52782 56194
rect 52782 56142 52834 56194
rect 52834 56142 52836 56194
rect 52780 56140 52836 56142
rect 49980 56082 50036 56084
rect 49980 56030 49982 56082
rect 49982 56030 50034 56082
rect 50034 56030 50036 56082
rect 49980 56028 50036 56030
rect 55132 56306 55188 56308
rect 55132 56254 55134 56306
rect 55134 56254 55186 56306
rect 55186 56254 55188 56306
rect 55132 56252 55188 56254
rect 55916 56252 55972 56308
rect 49868 55916 49924 55972
rect 50652 55970 50708 55972
rect 50652 55918 50654 55970
rect 50654 55918 50706 55970
rect 50706 55918 50708 55970
rect 50652 55916 50708 55918
rect 45500 53506 45556 53508
rect 45500 53454 45502 53506
rect 45502 53454 45554 53506
rect 45554 53454 45556 53506
rect 45500 53452 45556 53454
rect 46060 52220 46116 52276
rect 46060 50652 46116 50708
rect 44268 50034 44324 50036
rect 44268 49982 44270 50034
rect 44270 49982 44322 50034
rect 44322 49982 44324 50034
rect 44268 49980 44324 49982
rect 43372 46562 43428 46564
rect 43372 46510 43374 46562
rect 43374 46510 43426 46562
rect 43426 46510 43428 46562
rect 43372 46508 43428 46510
rect 43260 41074 43316 41076
rect 43260 41022 43262 41074
rect 43262 41022 43314 41074
rect 43314 41022 43316 41074
rect 43260 41020 43316 41022
rect 43148 40236 43204 40292
rect 43036 36764 43092 36820
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 51436 53564 51492 53620
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 57820 57708 57876 57764
rect 55580 52780 55636 52836
rect 58044 55356 58100 55412
rect 52668 52274 52724 52276
rect 52668 52222 52670 52274
rect 52670 52222 52722 52274
rect 52722 52222 52724 52274
rect 52668 52220 52724 52222
rect 51772 52162 51828 52164
rect 51772 52110 51774 52162
rect 51774 52110 51826 52162
rect 51826 52110 51828 52162
rect 51772 52108 51828 52110
rect 51548 51938 51604 51940
rect 51548 51886 51550 51938
rect 51550 51886 51602 51938
rect 51602 51886 51604 51938
rect 51548 51884 51604 51886
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 47068 50652 47124 50708
rect 46620 48524 46676 48580
rect 53452 52162 53508 52164
rect 53452 52110 53454 52162
rect 53454 52110 53506 52162
rect 53506 52110 53508 52162
rect 53452 52108 53508 52110
rect 52220 51884 52276 51940
rect 54124 52162 54180 52164
rect 54124 52110 54126 52162
rect 54126 52110 54178 52162
rect 54178 52110 54180 52162
rect 54124 52108 54180 52110
rect 51548 50540 51604 50596
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 47068 48300 47124 48356
rect 49084 48748 49140 48804
rect 47516 48636 47572 48692
rect 48188 48636 48244 48692
rect 47516 48188 47572 48244
rect 47852 48524 47908 48580
rect 48076 48354 48132 48356
rect 48076 48302 48078 48354
rect 48078 48302 48130 48354
rect 48130 48302 48132 48354
rect 48076 48300 48132 48302
rect 56252 52108 56308 52164
rect 55804 51324 55860 51380
rect 57260 50482 57316 50484
rect 57260 50430 57262 50482
rect 57262 50430 57314 50482
rect 57314 50430 57316 50482
rect 57260 50428 57316 50430
rect 58044 50482 58100 50484
rect 58044 50430 58046 50482
rect 58046 50430 58098 50482
rect 58098 50430 58100 50482
rect 58044 50428 58100 50430
rect 53116 48748 53172 48804
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 47740 46562 47796 46564
rect 47740 46510 47742 46562
rect 47742 46510 47794 46562
rect 47794 46510 47796 46562
rect 47740 46508 47796 46510
rect 48748 46562 48804 46564
rect 48748 46510 48750 46562
rect 48750 46510 48802 46562
rect 48802 46510 48804 46562
rect 48748 46508 48804 46510
rect 50092 46508 50148 46564
rect 47628 46450 47684 46452
rect 47628 46398 47630 46450
rect 47630 46398 47682 46450
rect 47682 46398 47684 46450
rect 47628 46396 47684 46398
rect 46508 45164 46564 45220
rect 43596 41244 43652 41300
rect 44156 41916 44212 41972
rect 43820 40962 43876 40964
rect 43820 40910 43822 40962
rect 43822 40910 43874 40962
rect 43874 40910 43876 40962
rect 43820 40908 43876 40910
rect 43372 40460 43428 40516
rect 45500 39340 45556 39396
rect 43708 38668 43764 38724
rect 43484 37436 43540 37492
rect 42140 36594 42196 36596
rect 42140 36542 42142 36594
rect 42142 36542 42194 36594
rect 42194 36542 42196 36594
rect 42140 36540 42196 36542
rect 41804 35308 41860 35364
rect 41020 30268 41076 30324
rect 41692 33068 41748 33124
rect 42700 34972 42756 35028
rect 42028 33458 42084 33460
rect 42028 33406 42030 33458
rect 42030 33406 42082 33458
rect 42082 33406 42084 33458
rect 42028 33404 42084 33406
rect 42476 33458 42532 33460
rect 42476 33406 42478 33458
rect 42478 33406 42530 33458
rect 42530 33406 42532 33458
rect 42476 33404 42532 33406
rect 41916 33346 41972 33348
rect 41916 33294 41918 33346
rect 41918 33294 41970 33346
rect 41970 33294 41972 33346
rect 41916 33292 41972 33294
rect 41356 31554 41412 31556
rect 41356 31502 41358 31554
rect 41358 31502 41410 31554
rect 41410 31502 41412 31554
rect 41356 31500 41412 31502
rect 41580 30882 41636 30884
rect 41580 30830 41582 30882
rect 41582 30830 41634 30882
rect 41634 30830 41636 30882
rect 41580 30828 41636 30830
rect 41244 28588 41300 28644
rect 41356 30156 41412 30212
rect 41692 28418 41748 28420
rect 41692 28366 41694 28418
rect 41694 28366 41746 28418
rect 41746 28366 41748 28418
rect 41692 28364 41748 28366
rect 41580 26402 41636 26404
rect 41580 26350 41582 26402
rect 41582 26350 41634 26402
rect 41634 26350 41636 26402
rect 41580 26348 41636 26350
rect 42140 31500 42196 31556
rect 42252 28364 42308 28420
rect 41916 26460 41972 26516
rect 42028 26908 42084 26964
rect 41132 17500 41188 17556
rect 40684 3164 40740 3220
rect 44604 38722 44660 38724
rect 44604 38670 44606 38722
rect 44606 38670 44658 38722
rect 44658 38670 44660 38722
rect 44604 38668 44660 38670
rect 43708 36428 43764 36484
rect 45500 39058 45556 39060
rect 45500 39006 45502 39058
rect 45502 39006 45554 39058
rect 45554 39006 45556 39058
rect 45500 39004 45556 39006
rect 45612 42028 45668 42084
rect 45388 38834 45444 38836
rect 45388 38782 45390 38834
rect 45390 38782 45442 38834
rect 45442 38782 45444 38834
rect 45388 38780 45444 38782
rect 44716 35756 44772 35812
rect 45164 36428 45220 36484
rect 45164 35644 45220 35700
rect 43148 34972 43204 35028
rect 44716 35026 44772 35028
rect 44716 34974 44718 35026
rect 44718 34974 44770 35026
rect 44770 34974 44772 35026
rect 44716 34972 44772 34974
rect 45164 34972 45220 35028
rect 45164 34354 45220 34356
rect 45164 34302 45166 34354
rect 45166 34302 45218 34354
rect 45218 34302 45220 34354
rect 45164 34300 45220 34302
rect 42700 32674 42756 32676
rect 42700 32622 42702 32674
rect 42702 32622 42754 32674
rect 42754 32622 42756 32674
rect 42700 32620 42756 32622
rect 42700 26514 42756 26516
rect 42700 26462 42702 26514
rect 42702 26462 42754 26514
rect 42754 26462 42756 26514
rect 42700 26460 42756 26462
rect 44268 3666 44324 3668
rect 44268 3614 44270 3666
rect 44270 3614 44322 3666
rect 44322 3614 44324 3666
rect 44268 3612 44324 3614
rect 42476 3500 42532 3556
rect 42364 3276 42420 3332
rect 48972 40908 49028 40964
rect 47516 39618 47572 39620
rect 47516 39566 47518 39618
rect 47518 39566 47570 39618
rect 47570 39566 47572 39618
rect 47516 39564 47572 39566
rect 47628 40236 47684 40292
rect 46732 39452 46788 39508
rect 47292 39506 47348 39508
rect 47292 39454 47294 39506
rect 47294 39454 47346 39506
rect 47346 39454 47348 39506
rect 47292 39452 47348 39454
rect 48188 40290 48244 40292
rect 48188 40238 48190 40290
rect 48190 40238 48242 40290
rect 48242 40238 48244 40290
rect 48188 40236 48244 40238
rect 47628 39452 47684 39508
rect 47852 39452 47908 39508
rect 48748 39506 48804 39508
rect 48748 39454 48750 39506
rect 48750 39454 48802 39506
rect 48802 39454 48804 39506
rect 48748 39452 48804 39454
rect 46620 39058 46676 39060
rect 46620 39006 46622 39058
rect 46622 39006 46674 39058
rect 46674 39006 46676 39058
rect 46620 39004 46676 39006
rect 45948 38834 46004 38836
rect 45948 38782 45950 38834
rect 45950 38782 46002 38834
rect 46002 38782 46004 38834
rect 45948 38780 46004 38782
rect 49644 39452 49700 39508
rect 48524 38780 48580 38836
rect 45724 38722 45780 38724
rect 45724 38670 45726 38722
rect 45726 38670 45778 38722
rect 45778 38670 45780 38722
rect 45724 38668 45780 38670
rect 46060 36876 46116 36932
rect 45948 35922 46004 35924
rect 45948 35870 45950 35922
rect 45950 35870 46002 35922
rect 46002 35870 46004 35922
rect 45948 35868 46004 35870
rect 45836 35810 45892 35812
rect 45836 35758 45838 35810
rect 45838 35758 45890 35810
rect 45890 35758 45892 35810
rect 45836 35756 45892 35758
rect 46060 35756 46116 35812
rect 49980 36988 50036 37044
rect 47292 35810 47348 35812
rect 47292 35758 47294 35810
rect 47294 35758 47346 35810
rect 47346 35758 47348 35810
rect 47292 35756 47348 35758
rect 46284 35698 46340 35700
rect 46284 35646 46286 35698
rect 46286 35646 46338 35698
rect 46338 35646 46340 35698
rect 46284 35644 46340 35646
rect 46508 35698 46564 35700
rect 46508 35646 46510 35698
rect 46510 35646 46562 35698
rect 46562 35646 46564 35698
rect 46508 35644 46564 35646
rect 45836 34354 45892 34356
rect 45836 34302 45838 34354
rect 45838 34302 45890 34354
rect 45890 34302 45892 34354
rect 45836 34300 45892 34302
rect 45948 34412 46004 34468
rect 49420 35644 49476 35700
rect 49308 35196 49364 35252
rect 49532 35196 49588 35252
rect 46732 34412 46788 34468
rect 49980 35196 50036 35252
rect 52892 46060 52948 46116
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50876 40572 50932 40628
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50988 36988 51044 37044
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50092 35698 50148 35700
rect 50092 35646 50094 35698
rect 50094 35646 50146 35698
rect 50146 35646 50148 35698
rect 50092 35644 50148 35646
rect 50876 35698 50932 35700
rect 50876 35646 50878 35698
rect 50878 35646 50930 35698
rect 50930 35646 50932 35698
rect 50876 35644 50932 35646
rect 50092 33122 50148 33124
rect 50092 33070 50094 33122
rect 50094 33070 50146 33122
rect 50146 33070 50148 33122
rect 50092 33068 50148 33070
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50316 33068 50372 33124
rect 50540 33122 50596 33124
rect 50540 33070 50542 33122
rect 50542 33070 50594 33122
rect 50594 33070 50596 33122
rect 50540 33068 50596 33070
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 51884 35698 51940 35700
rect 51884 35646 51886 35698
rect 51886 35646 51938 35698
rect 51938 35646 51940 35698
rect 51884 35644 51940 35646
rect 51324 35420 51380 35476
rect 57260 43820 57316 43876
rect 57596 42812 57652 42868
rect 58044 43820 58100 43876
rect 57260 41074 57316 41076
rect 57260 41022 57262 41074
rect 57262 41022 57314 41074
rect 57314 41022 57316 41074
rect 57260 41020 57316 41022
rect 58044 41074 58100 41076
rect 58044 41022 58046 41074
rect 58046 41022 58098 41074
rect 58098 41022 58100 41074
rect 58044 41020 58100 41022
rect 57708 40348 57764 40404
rect 57596 37884 57652 37940
rect 57260 37826 57316 37828
rect 57260 37774 57262 37826
rect 57262 37774 57314 37826
rect 57314 37774 57316 37826
rect 57260 37772 57316 37774
rect 58044 37772 58100 37828
rect 57708 37436 57764 37492
rect 52892 34972 52948 35028
rect 56252 35026 56308 35028
rect 56252 34974 56254 35026
rect 56254 34974 56306 35026
rect 56306 34974 56308 35026
rect 56252 34972 56308 34974
rect 56812 34972 56868 35028
rect 57820 35026 57876 35028
rect 57820 34974 57822 35026
rect 57822 34974 57874 35026
rect 57874 34974 57876 35026
rect 57820 34972 57876 34974
rect 57708 33068 57764 33124
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 46732 23212 46788 23268
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 46508 20636 46564 20692
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 57484 31164 57540 31220
rect 56252 27692 56308 27748
rect 57260 20300 57316 20356
rect 57260 17442 57316 17444
rect 57260 17390 57262 17442
rect 57262 17390 57314 17442
rect 57314 17390 57316 17442
rect 57260 17388 57316 17390
rect 51324 14588 51380 14644
rect 56364 14642 56420 14644
rect 56364 14590 56366 14642
rect 56366 14590 56418 14642
rect 56418 14590 56420 14642
rect 56364 14588 56420 14590
rect 56812 14588 56868 14644
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 56364 11170 56420 11172
rect 56364 11118 56366 11170
rect 56366 11118 56418 11170
rect 56418 11118 56420 11170
rect 56364 11116 56420 11118
rect 56812 11116 56868 11172
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 57596 30828 57652 30884
rect 58044 31554 58100 31556
rect 58044 31502 58046 31554
rect 58046 31502 58098 31554
rect 58098 31502 58100 31554
rect 58044 31500 58100 31502
rect 58156 28812 58212 28868
rect 57820 25618 57876 25620
rect 57820 25566 57822 25618
rect 57822 25566 57874 25618
rect 57874 25566 57876 25618
rect 57820 25564 57876 25566
rect 57708 23266 57764 23268
rect 57708 23214 57710 23266
rect 57710 23214 57762 23266
rect 57762 23214 57764 23266
rect 57708 23212 57764 23214
rect 58044 22988 58100 23044
rect 57708 20690 57764 20692
rect 57708 20638 57710 20690
rect 57710 20638 57762 20690
rect 57762 20638 57764 20690
rect 57708 20636 57764 20638
rect 58044 20300 58100 20356
rect 57708 17554 57764 17556
rect 57708 17502 57710 17554
rect 57710 17502 57762 17554
rect 57762 17502 57764 17554
rect 57708 17500 57764 17502
rect 57708 14252 57764 14308
rect 57708 10892 57764 10948
rect 57260 8034 57316 8036
rect 57260 7982 57262 8034
rect 57262 7982 57314 8034
rect 57314 7982 57316 8034
rect 57260 7980 57316 7982
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 57260 5010 57316 5012
rect 57260 4958 57262 5010
rect 57262 4958 57314 5010
rect 57314 4958 57316 5010
rect 57260 4956 57316 4958
rect 57708 8146 57764 8148
rect 57708 8094 57710 8146
rect 57710 8094 57762 8146
rect 57762 8094 57764 8146
rect 57708 8092 57764 8094
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 58044 17388 58100 17444
rect 58044 16940 58100 16996
rect 58044 8146 58100 8148
rect 58044 8094 58046 8146
rect 58046 8094 58098 8146
rect 58098 8094 58100 8146
rect 58044 8092 58100 8094
rect 58044 5180 58100 5236
rect 58044 5010 58100 5012
rect 58044 4958 58046 5010
rect 58046 4958 58098 5010
rect 58098 4958 58100 5010
rect 58044 4956 58100 4958
rect 56812 4226 56868 4228
rect 56812 4174 56814 4226
rect 56814 4174 56866 4226
rect 56866 4174 56868 4226
rect 56812 4172 56868 4174
rect 58044 4172 58100 4228
rect 45612 3612 45668 3668
rect 56028 3554 56084 3556
rect 56028 3502 56030 3554
rect 56030 3502 56082 3554
rect 56082 3502 56084 3554
rect 56028 3500 56084 3502
rect 56700 3554 56756 3556
rect 56700 3502 56702 3554
rect 56702 3502 56754 3554
rect 56754 3502 56756 3554
rect 56700 3500 56756 3502
rect 48188 3442 48244 3444
rect 48188 3390 48190 3442
rect 48190 3390 48242 3442
rect 48242 3390 48244 3442
rect 48188 3388 48244 3390
rect 49196 3442 49252 3444
rect 49196 3390 49198 3442
rect 49198 3390 49250 3442
rect 49250 3390 49252 3442
rect 49196 3388 49252 3390
rect 50428 3388 50484 3444
rect 48860 3164 48916 3220
rect 50988 3442 51044 3444
rect 50988 3390 50990 3442
rect 50990 3390 51042 3442
rect 51042 3390 51044 3442
rect 50988 3388 51044 3390
rect 56588 3388 56644 3444
rect 50652 3330 50708 3332
rect 50652 3278 50654 3330
rect 50654 3278 50706 3330
rect 50706 3278 50708 3330
rect 50652 3276 50708 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 57596 3442 57652 3444
rect 57596 3390 57598 3442
rect 57598 3390 57650 3442
rect 57650 3390 57652 3442
rect 57596 3388 57652 3390
rect 58044 2828 58100 2884
<< metal3 >>
rect 200 59080 800 59304
rect 59200 58436 59800 58632
rect 59164 58408 59800 58436
rect 59164 58380 59304 58408
rect 59164 58324 59220 58380
rect 59164 58268 59332 58324
rect 59276 57764 59332 58268
rect 57810 57708 57820 57764
rect 57876 57708 59332 57764
rect 200 56420 800 56616
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 200 56392 1820 56420
rect 728 56364 1820 56392
rect 1876 56364 1886 56420
rect 55122 56252 55132 56308
rect 55188 56252 55916 56308
rect 55972 56252 55982 56308
rect 4834 56140 4844 56196
rect 4900 56140 6076 56196
rect 6132 56140 6142 56196
rect 28354 56140 28364 56196
rect 28420 56140 31836 56196
rect 31892 56140 31902 56196
rect 38210 56140 38220 56196
rect 38276 56140 39788 56196
rect 39844 56140 39854 56196
rect 41122 56140 41132 56196
rect 41188 56140 42140 56196
rect 42196 56140 42206 56196
rect 44930 56140 44940 56196
rect 44996 56140 52780 56196
rect 52836 56140 52846 56196
rect 25330 56028 25340 56084
rect 25396 56028 26796 56084
rect 26852 56028 26862 56084
rect 31490 56028 31500 56084
rect 31556 56028 32060 56084
rect 32116 56028 32126 56084
rect 42578 56028 42588 56084
rect 42644 56028 49532 56084
rect 49588 56028 49980 56084
rect 50036 56028 50046 56084
rect 3490 55916 3500 55972
rect 3556 55916 4060 55972
rect 4116 55916 7644 55972
rect 7700 55916 7710 55972
rect 18722 55916 18732 55972
rect 18788 55916 20636 55972
rect 20692 55916 22764 55972
rect 22820 55916 22830 55972
rect 49858 55916 49868 55972
rect 49924 55916 50652 55972
rect 50708 55916 50718 55972
rect 18834 55804 18844 55860
rect 18900 55804 22652 55860
rect 22708 55804 24108 55860
rect 24164 55804 24174 55860
rect 59200 55748 59800 55944
rect 59164 55720 59800 55748
rect 59164 55692 59304 55720
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 59164 55636 59220 55692
rect 59164 55580 59332 55636
rect 59276 55412 59332 55580
rect 40338 55356 40348 55412
rect 40404 55356 41244 55412
rect 41300 55356 41310 55412
rect 58034 55356 58044 55412
rect 58100 55356 59332 55412
rect 17938 55132 17948 55188
rect 18004 55132 28588 55188
rect 28644 55132 29260 55188
rect 29316 55132 29326 55188
rect 8306 55020 8316 55076
rect 8372 54852 8428 55076
rect 10770 55020 10780 55076
rect 10836 55020 12348 55076
rect 12404 55020 15260 55076
rect 15316 55020 15326 55076
rect 18722 55020 18732 55076
rect 18788 55020 20860 55076
rect 20916 55020 20926 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 8372 54796 11452 54852
rect 11508 54796 11518 54852
rect 20178 54684 20188 54740
rect 20244 54684 38444 54740
rect 38500 54684 38510 54740
rect 19282 54572 19292 54628
rect 19348 54572 28476 54628
rect 28532 54572 40348 54628
rect 40404 54572 40414 54628
rect 16258 54460 16268 54516
rect 16324 54460 19404 54516
rect 19460 54460 20300 54516
rect 20356 54460 20366 54516
rect 20738 54348 20748 54404
rect 20804 54348 24220 54404
rect 24276 54348 35980 54404
rect 36036 54348 36046 54404
rect 11442 54236 11452 54292
rect 11508 54236 28700 54292
rect 28756 54236 28766 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 20850 53900 20860 53956
rect 20916 53900 30268 53956
rect 30324 53900 30334 53956
rect 2034 53788 2044 53844
rect 2100 53788 3724 53844
rect 3780 53788 3790 53844
rect 39218 53788 39228 53844
rect 39284 53788 42364 53844
rect 42420 53788 42430 53844
rect 9090 53676 9100 53732
rect 9156 53676 12460 53732
rect 12516 53676 12526 53732
rect 13794 53676 13804 53732
rect 13860 53676 14812 53732
rect 14868 53676 14878 53732
rect 17378 53676 17388 53732
rect 17444 53676 18732 53732
rect 18788 53676 32508 53732
rect 32564 53676 32574 53732
rect 12114 53564 12124 53620
rect 12180 53564 18844 53620
rect 18900 53564 18910 53620
rect 23202 53564 23212 53620
rect 23268 53564 27356 53620
rect 27412 53564 27422 53620
rect 27794 53564 27804 53620
rect 27860 53564 28812 53620
rect 28868 53564 29148 53620
rect 29204 53564 29214 53620
rect 29474 53564 29484 53620
rect 29540 53564 30380 53620
rect 30436 53564 30716 53620
rect 30772 53564 31052 53620
rect 31108 53564 31118 53620
rect 42130 53564 42140 53620
rect 42196 53564 42812 53620
rect 42868 53564 51436 53620
rect 51492 53564 51502 53620
rect 29148 53508 29204 53564
rect 11890 53452 11900 53508
rect 11956 53452 12684 53508
rect 12740 53452 12750 53508
rect 29148 53452 30492 53508
rect 30548 53452 30558 53508
rect 39106 53452 39116 53508
rect 39172 53452 39564 53508
rect 39620 53452 40012 53508
rect 40068 53452 40684 53508
rect 40740 53452 40750 53508
rect 41682 53452 41692 53508
rect 41748 53452 45500 53508
rect 45556 53452 45566 53508
rect 40786 53340 40796 53396
rect 40852 53340 41468 53396
rect 41524 53340 41534 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 200 53172 800 53256
rect 23212 53228 29708 53284
rect 29764 53228 29774 53284
rect 23212 53172 23268 53228
rect 200 53116 1820 53172
rect 1876 53116 1886 53172
rect 11554 53116 11564 53172
rect 11620 53116 12348 53172
rect 12404 53116 23268 53172
rect 23426 53116 23436 53172
rect 23492 53116 29036 53172
rect 29092 53116 29102 53172
rect 200 53032 800 53116
rect 2258 53004 2268 53060
rect 2324 53004 3724 53060
rect 3780 53004 3790 53060
rect 6178 53004 6188 53060
rect 6244 53004 10556 53060
rect 10612 53004 10622 53060
rect 14130 53004 14140 53060
rect 14196 53004 18620 53060
rect 18676 53004 20188 53060
rect 28018 53004 28028 53060
rect 28084 53004 42700 53060
rect 42756 53004 43372 53060
rect 43428 53004 43438 53060
rect 20132 52948 20188 53004
rect 8194 52892 8204 52948
rect 8260 52892 8652 52948
rect 8708 52892 9100 52948
rect 9156 52892 9660 52948
rect 9716 52892 9726 52948
rect 16482 52892 16492 52948
rect 16548 52892 18172 52948
rect 18228 52892 18238 52948
rect 20132 52892 30940 52948
rect 30996 52892 31006 52948
rect 3938 52780 3948 52836
rect 4004 52780 4508 52836
rect 4564 52780 4574 52836
rect 8530 52780 8540 52836
rect 8596 52780 10220 52836
rect 10276 52780 10286 52836
rect 19506 52780 19516 52836
rect 19572 52780 19964 52836
rect 20020 52780 20524 52836
rect 20580 52780 20590 52836
rect 27346 52780 27356 52836
rect 27412 52780 29820 52836
rect 29876 52780 29886 52836
rect 43586 52780 43596 52836
rect 43652 52780 44044 52836
rect 44100 52780 55580 52836
rect 55636 52780 55646 52836
rect 24098 52668 24108 52724
rect 24164 52668 25340 52724
rect 25396 52668 25900 52724
rect 25956 52668 25966 52724
rect 10546 52556 10556 52612
rect 10612 52556 31388 52612
rect 31444 52556 31454 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 59200 52360 59800 52584
rect 10210 52220 10220 52276
rect 10276 52220 11900 52276
rect 11956 52220 15148 52276
rect 15204 52220 15214 52276
rect 16930 52220 16940 52276
rect 16996 52220 18956 52276
rect 19012 52220 21532 52276
rect 21588 52220 21598 52276
rect 28466 52220 28476 52276
rect 28532 52220 29148 52276
rect 29204 52220 29484 52276
rect 29540 52220 29550 52276
rect 30034 52220 30044 52276
rect 30100 52220 32620 52276
rect 32676 52220 32686 52276
rect 46050 52220 46060 52276
rect 46116 52220 52668 52276
rect 52724 52220 54180 52276
rect 54124 52164 54180 52220
rect 9650 52108 9660 52164
rect 9716 52108 10892 52164
rect 10948 52108 11452 52164
rect 11508 52108 12684 52164
rect 12740 52108 12750 52164
rect 14466 52108 14476 52164
rect 14532 52108 15036 52164
rect 15092 52108 15820 52164
rect 15876 52108 16492 52164
rect 16548 52108 17052 52164
rect 17108 52108 17612 52164
rect 17668 52108 18284 52164
rect 18340 52108 18350 52164
rect 22642 52108 22652 52164
rect 22708 52108 28364 52164
rect 28420 52108 28430 52164
rect 30706 52108 30716 52164
rect 30772 52108 35532 52164
rect 35588 52108 35598 52164
rect 39890 52108 39900 52164
rect 39956 52108 40796 52164
rect 40852 52108 40862 52164
rect 51762 52108 51772 52164
rect 51828 52108 53452 52164
rect 53508 52108 53518 52164
rect 54114 52108 54124 52164
rect 54180 52108 56252 52164
rect 56308 52108 56318 52164
rect 21074 51996 21084 52052
rect 21140 51996 24556 52052
rect 24612 51996 25228 52052
rect 25284 51996 25294 52052
rect 7970 51884 7980 51940
rect 8036 51884 11116 51940
rect 11172 51884 11182 51940
rect 51538 51884 51548 51940
rect 51604 51884 52220 51940
rect 52276 51884 52286 51940
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 19730 51548 19740 51604
rect 19796 51548 41244 51604
rect 41300 51548 41310 51604
rect 2146 51436 2156 51492
rect 2212 51436 4620 51492
rect 4676 51436 4686 51492
rect 18050 51436 18060 51492
rect 18116 51436 18732 51492
rect 18788 51436 31052 51492
rect 31108 51436 31118 51492
rect 40226 51436 40236 51492
rect 40292 51436 41468 51492
rect 41524 51436 41534 51492
rect 11106 51324 11116 51380
rect 11172 51324 30380 51380
rect 30436 51324 30446 51380
rect 39900 51324 40684 51380
rect 40740 51324 40750 51380
rect 42466 51324 42476 51380
rect 42532 51324 43484 51380
rect 43540 51324 55804 51380
rect 55860 51324 55870 51380
rect 39900 51268 39956 51324
rect 37538 51212 37548 51268
rect 37604 51212 38556 51268
rect 38612 51212 39900 51268
rect 39956 51212 39966 51268
rect 3378 51100 3388 51156
rect 3444 51100 4732 51156
rect 4788 51100 4798 51156
rect 29810 51100 29820 51156
rect 29876 51100 42140 51156
rect 42196 51100 43148 51156
rect 43204 51100 43214 51156
rect 39442 50988 39452 51044
rect 39508 50988 40236 51044
rect 40292 50988 40302 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 22082 50876 22092 50932
rect 22148 50876 27244 50932
rect 27300 50876 27310 50932
rect 10322 50764 10332 50820
rect 10388 50764 40012 50820
rect 40068 50764 40078 50820
rect 40450 50764 40460 50820
rect 40516 50764 43036 50820
rect 43092 50764 43102 50820
rect 18610 50652 18620 50708
rect 18676 50652 46060 50708
rect 46116 50652 47068 50708
rect 47124 50652 47134 50708
rect 200 50484 800 50568
rect 15586 50540 15596 50596
rect 15652 50540 19740 50596
rect 19796 50540 19806 50596
rect 43652 50540 51548 50596
rect 51604 50540 51614 50596
rect 43652 50484 43708 50540
rect 200 50428 1820 50484
rect 1876 50428 1886 50484
rect 8642 50428 8652 50484
rect 8708 50428 11228 50484
rect 11284 50428 12684 50484
rect 12740 50428 12750 50484
rect 36754 50428 36764 50484
rect 36820 50428 39452 50484
rect 39508 50428 39518 50484
rect 40226 50428 40236 50484
rect 40292 50428 40908 50484
rect 40964 50428 43708 50484
rect 57250 50428 57260 50484
rect 57316 50428 58044 50484
rect 58100 50428 59332 50484
rect 200 50344 800 50428
rect 3938 50316 3948 50372
rect 4004 50316 5180 50372
rect 5236 50316 5246 50372
rect 19170 50316 19180 50372
rect 19236 50316 19516 50372
rect 19572 50316 19582 50372
rect 20178 50316 20188 50372
rect 20244 50316 23660 50372
rect 23716 50316 23726 50372
rect 19058 50204 19068 50260
rect 19124 50204 19134 50260
rect 19068 50036 19124 50204
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 59276 50036 59332 50428
rect 19068 49980 22204 50036
rect 22260 49980 22270 50036
rect 43586 49980 43596 50036
rect 43652 49980 44268 50036
rect 44324 49980 44334 50036
rect 59164 49980 59332 50036
rect 59164 49924 59220 49980
rect 10994 49868 11004 49924
rect 11060 49868 11452 49924
rect 11508 49868 12236 49924
rect 12292 49868 12302 49924
rect 15250 49868 15260 49924
rect 15316 49868 30380 49924
rect 30436 49868 30446 49924
rect 32162 49868 32172 49924
rect 32228 49868 32396 49924
rect 32452 49868 32620 49924
rect 32676 49868 35868 49924
rect 35924 49868 35934 49924
rect 59164 49896 59304 49924
rect 59164 49868 59800 49896
rect 15026 49756 15036 49812
rect 15092 49756 15596 49812
rect 15652 49756 15662 49812
rect 18498 49756 18508 49812
rect 18564 49756 18956 49812
rect 19012 49756 19180 49812
rect 19236 49756 19246 49812
rect 23650 49756 23660 49812
rect 23716 49756 37772 49812
rect 37828 49756 37838 49812
rect 19618 49644 19628 49700
rect 19684 49644 23100 49700
rect 23156 49644 28364 49700
rect 28420 49644 28430 49700
rect 31490 49644 31500 49700
rect 31556 49644 32172 49700
rect 32228 49644 32238 49700
rect 59200 49672 59800 49868
rect 11106 49532 11116 49588
rect 11172 49532 11900 49588
rect 11956 49532 32060 49588
rect 32116 49532 32126 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 32498 49084 32508 49140
rect 32564 49084 35868 49140
rect 35924 49084 35934 49140
rect 4050 48972 4060 49028
rect 4116 48972 4956 49028
rect 5012 48972 5022 49028
rect 8372 48860 10556 48916
rect 10612 48860 31836 48916
rect 31892 48860 31902 48916
rect 8372 48804 8428 48860
rect 2146 48748 2156 48804
rect 2212 48748 3724 48804
rect 3780 48748 3790 48804
rect 4498 48748 4508 48804
rect 4564 48748 5180 48804
rect 5236 48748 6580 48804
rect 7410 48748 7420 48804
rect 7476 48748 8428 48804
rect 9762 48748 9772 48804
rect 9828 48748 11340 48804
rect 11396 48748 12796 48804
rect 12852 48748 12862 48804
rect 15586 48748 15596 48804
rect 15652 48748 18396 48804
rect 18452 48748 20524 48804
rect 20580 48748 21532 48804
rect 21588 48748 21598 48804
rect 22194 48748 22204 48804
rect 22260 48748 29596 48804
rect 29652 48748 29662 48804
rect 36418 48748 36428 48804
rect 36484 48748 36988 48804
rect 37044 48748 37436 48804
rect 37492 48748 37502 48804
rect 48748 48748 49084 48804
rect 49140 48748 53116 48804
rect 53172 48748 53182 48804
rect 6524 48580 6580 48748
rect 48748 48692 48804 48748
rect 13122 48636 13132 48692
rect 13188 48636 13804 48692
rect 13860 48636 13870 48692
rect 33842 48636 33852 48692
rect 33908 48636 39004 48692
rect 39060 48636 43708 48692
rect 47506 48636 47516 48692
rect 47572 48636 48188 48692
rect 48244 48636 48804 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 43652 48580 43708 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 6514 48524 6524 48580
rect 6580 48524 6590 48580
rect 43652 48524 46620 48580
rect 46676 48524 47852 48580
rect 47908 48524 47918 48580
rect 11442 48412 11452 48468
rect 11508 48412 12124 48468
rect 12180 48412 31388 48468
rect 31444 48412 31454 48468
rect 3938 48300 3948 48356
rect 4004 48300 4508 48356
rect 4564 48300 4574 48356
rect 18162 48300 18172 48356
rect 18228 48300 36764 48356
rect 36820 48300 36830 48356
rect 47058 48300 47068 48356
rect 47124 48300 48076 48356
rect 48132 48300 48142 48356
rect 26562 48188 26572 48244
rect 26628 48188 47516 48244
rect 47572 48188 47582 48244
rect 23202 48076 23212 48132
rect 23268 48076 37996 48132
rect 38052 48076 38556 48132
rect 38612 48076 42476 48132
rect 42532 48076 42542 48132
rect 15138 47964 15148 48020
rect 15204 47964 43036 48020
rect 43092 47964 43102 48020
rect 728 47880 2044 47908
rect 200 47852 2044 47880
rect 2100 47852 2110 47908
rect 200 47656 800 47852
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 5394 47516 5404 47572
rect 5460 47516 5852 47572
rect 5908 47516 8428 47572
rect 14018 47516 14028 47572
rect 14084 47516 19404 47572
rect 19460 47516 19470 47572
rect 26786 47516 26796 47572
rect 26852 47516 27356 47572
rect 27412 47516 27422 47572
rect 8372 47460 8428 47516
rect 8372 47404 31612 47460
rect 31668 47404 31678 47460
rect 3826 47292 3836 47348
rect 3892 47292 4844 47348
rect 4900 47292 4910 47348
rect 23426 47180 23436 47236
rect 23492 47180 27916 47236
rect 27972 47180 27982 47236
rect 2034 47068 2044 47124
rect 2100 47068 3724 47124
rect 3780 47068 3790 47124
rect 23314 47068 23324 47124
rect 23380 47068 28588 47124
rect 28644 47068 28654 47124
rect 38322 47068 38332 47124
rect 38388 47068 40124 47124
rect 40180 47068 40190 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 28018 46956 28028 47012
rect 28084 46956 28252 47012
rect 28308 46956 28700 47012
rect 28756 46956 29484 47012
rect 29540 46956 29932 47012
rect 29988 46956 31724 47012
rect 31780 46956 31790 47012
rect 59200 46984 59800 47208
rect 3164 46620 3724 46676
rect 3780 46620 3790 46676
rect 41794 46620 41804 46676
rect 41860 46620 42924 46676
rect 42980 46620 42990 46676
rect 3164 46564 3220 46620
rect 2482 46508 2492 46564
rect 2548 46508 3164 46564
rect 3220 46508 3230 46564
rect 9090 46508 9100 46564
rect 9156 46508 12348 46564
rect 12404 46508 12414 46564
rect 16930 46508 16940 46564
rect 16996 46508 20076 46564
rect 20132 46508 29372 46564
rect 29428 46508 29438 46564
rect 32946 46508 32956 46564
rect 33012 46508 33740 46564
rect 33796 46508 33806 46564
rect 42354 46508 42364 46564
rect 42420 46508 43372 46564
rect 43428 46508 43438 46564
rect 47730 46508 47740 46564
rect 47796 46508 48748 46564
rect 48804 46508 50092 46564
rect 50148 46508 50158 46564
rect 21074 46396 21084 46452
rect 21140 46396 23548 46452
rect 23604 46396 24556 46452
rect 24612 46396 24622 46452
rect 41570 46396 41580 46452
rect 41636 46396 47628 46452
rect 47684 46396 47694 46452
rect 24070 46284 24108 46340
rect 24164 46284 24174 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 24098 46060 24108 46116
rect 24164 46060 52892 46116
rect 52948 46060 52958 46116
rect 10658 45948 10668 46004
rect 10724 45948 11228 46004
rect 11284 45948 12572 46004
rect 12628 45948 12638 46004
rect 13916 45948 21868 46004
rect 21924 45948 21934 46004
rect 13916 45892 13972 45948
rect 10098 45836 10108 45892
rect 10164 45836 11676 45892
rect 11732 45836 13972 45892
rect 19170 45836 19180 45892
rect 19236 45836 20860 45892
rect 20916 45836 20926 45892
rect 30706 45836 30716 45892
rect 30772 45836 31164 45892
rect 31220 45836 31230 45892
rect 35634 45836 35644 45892
rect 35700 45836 36652 45892
rect 36708 45836 36718 45892
rect 37090 45836 37100 45892
rect 37156 45836 37996 45892
rect 38052 45836 38062 45892
rect 15092 45724 16156 45780
rect 16212 45724 32620 45780
rect 32676 45724 32686 45780
rect 34066 45724 34076 45780
rect 34132 45724 34524 45780
rect 34580 45724 36988 45780
rect 37044 45724 41020 45780
rect 41076 45724 41086 45780
rect 15092 45668 15148 45724
rect 3266 45612 3276 45668
rect 3332 45612 15148 45668
rect 19394 45612 19404 45668
rect 19460 45612 19740 45668
rect 19796 45612 19806 45668
rect 30940 45612 37884 45668
rect 37940 45612 39004 45668
rect 39060 45612 39070 45668
rect 23492 45500 30716 45556
rect 30772 45500 30782 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 23492 45332 23548 45500
rect 30940 45444 30996 45612
rect 31154 45500 31164 45556
rect 31220 45500 35980 45556
rect 36036 45500 36046 45556
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 30930 45388 30940 45444
rect 30996 45388 31006 45444
rect 31490 45388 31500 45444
rect 31556 45388 31724 45444
rect 31780 45388 31790 45444
rect 40786 45388 40796 45444
rect 40852 45388 41916 45444
rect 41972 45388 43148 45444
rect 43204 45388 43214 45444
rect 7746 45276 7756 45332
rect 7812 45276 10780 45332
rect 10836 45276 10846 45332
rect 17378 45276 17388 45332
rect 17444 45276 23548 45332
rect 27570 45276 27580 45332
rect 27636 45276 29260 45332
rect 29316 45276 29326 45332
rect 29922 45276 29932 45332
rect 29988 45276 30716 45332
rect 30772 45276 33628 45332
rect 33684 45276 33694 45332
rect 38546 45276 38556 45332
rect 38612 45276 39900 45332
rect 39956 45276 39966 45332
rect 6178 45164 6188 45220
rect 6244 45164 9884 45220
rect 9940 45164 9950 45220
rect 24882 45164 24892 45220
rect 24948 45164 28588 45220
rect 28644 45164 28654 45220
rect 30258 45164 30268 45220
rect 30324 45164 30604 45220
rect 30660 45164 31164 45220
rect 31220 45164 31948 45220
rect 32004 45164 32172 45220
rect 32228 45164 32620 45220
rect 32676 45164 32686 45220
rect 37314 45164 37324 45220
rect 37380 45164 38220 45220
rect 38276 45164 46508 45220
rect 46564 45164 46574 45220
rect 8530 45052 8540 45108
rect 8596 45052 9436 45108
rect 9492 45052 11228 45108
rect 11284 45052 11294 45108
rect 20738 45052 20748 45108
rect 20804 45052 24332 45108
rect 24388 45052 24398 45108
rect 28690 45052 28700 45108
rect 28756 45052 29708 45108
rect 29764 45052 29774 45108
rect 30370 45052 30380 45108
rect 30436 45052 30828 45108
rect 30884 45052 30894 45108
rect 27906 44940 27916 44996
rect 27972 44940 29932 44996
rect 29988 44940 30156 44996
rect 30212 44940 30222 44996
rect 36642 44940 36652 44996
rect 36708 44940 36988 44996
rect 37044 44940 37772 44996
rect 37828 44940 37838 44996
rect 40002 44940 40012 44996
rect 40068 44940 41244 44996
rect 41300 44940 41580 44996
rect 41636 44940 41646 44996
rect 10770 44828 10780 44884
rect 10836 44828 31388 44884
rect 31444 44828 31454 44884
rect 9762 44716 9772 44772
rect 9828 44716 32060 44772
rect 32116 44716 32126 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 200 44436 800 44520
rect 29586 44492 29596 44548
rect 29652 44492 30156 44548
rect 30212 44492 30222 44548
rect 200 44380 1820 44436
rect 1876 44380 1886 44436
rect 28802 44380 28812 44436
rect 28868 44380 30268 44436
rect 30324 44380 30334 44436
rect 31602 44380 31612 44436
rect 31668 44380 33516 44436
rect 33572 44380 33582 44436
rect 200 44296 800 44380
rect 10546 44268 10556 44324
rect 10612 44268 12124 44324
rect 12180 44268 12190 44324
rect 17714 44268 17724 44324
rect 17780 44268 31052 44324
rect 31108 44268 31118 44324
rect 33618 44268 33628 44324
rect 33684 44268 34076 44324
rect 34132 44268 34142 44324
rect 17938 44156 17948 44212
rect 18004 44156 19292 44212
rect 19348 44156 33964 44212
rect 34020 44156 34030 44212
rect 8082 44044 8092 44100
rect 8148 44044 14364 44100
rect 14420 44044 15372 44100
rect 15428 44044 15438 44100
rect 18834 44044 18844 44100
rect 18900 44044 19628 44100
rect 19684 44044 19694 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 57250 43820 57260 43876
rect 57316 43820 58044 43876
rect 58100 43848 59304 43876
rect 58100 43820 59800 43848
rect 6178 43708 6188 43764
rect 6244 43708 9772 43764
rect 9828 43708 9838 43764
rect 16146 43708 16156 43764
rect 16212 43708 17724 43764
rect 17780 43708 17790 43764
rect 23426 43708 23436 43764
rect 23492 43708 24892 43764
rect 24948 43708 24958 43764
rect 9538 43596 9548 43652
rect 9604 43596 10220 43652
rect 10276 43596 15148 43652
rect 20962 43596 20972 43652
rect 21028 43596 24332 43652
rect 24388 43596 30044 43652
rect 30100 43596 30110 43652
rect 31266 43596 31276 43652
rect 31332 43596 31612 43652
rect 31668 43596 32060 43652
rect 32116 43596 33068 43652
rect 33124 43596 33134 43652
rect 34178 43596 34188 43652
rect 34244 43596 36876 43652
rect 36932 43596 36942 43652
rect 59200 43624 59800 43820
rect 15092 43540 15148 43596
rect 12674 43484 12684 43540
rect 12740 43484 13580 43540
rect 13636 43484 13646 43540
rect 15092 43484 34300 43540
rect 34356 43484 34366 43540
rect 36642 43484 36652 43540
rect 36708 43484 37660 43540
rect 37716 43484 37726 43540
rect 8866 43372 8876 43428
rect 8932 43372 9660 43428
rect 9716 43372 10108 43428
rect 10164 43372 10668 43428
rect 10724 43372 11116 43428
rect 11172 43372 11676 43428
rect 11732 43372 12124 43428
rect 12180 43372 12908 43428
rect 12964 43372 12974 43428
rect 32610 43372 32620 43428
rect 32676 43372 34188 43428
rect 34244 43372 34254 43428
rect 35970 43372 35980 43428
rect 36036 43372 37100 43428
rect 37156 43372 37996 43428
rect 38052 43372 38062 43428
rect 8194 43260 8204 43316
rect 8260 43260 11340 43316
rect 11396 43260 11406 43316
rect 23986 43260 23996 43316
rect 24052 43260 32396 43316
rect 32452 43260 32956 43316
rect 33012 43260 33022 43316
rect 35074 43260 35084 43316
rect 35140 43260 37324 43316
rect 37380 43260 37390 43316
rect 8530 43148 8540 43204
rect 8596 43148 10780 43204
rect 10836 43148 15820 43204
rect 15876 43148 15886 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 9874 43036 9884 43092
rect 9940 43036 31500 43092
rect 31556 43036 31566 43092
rect 11330 42924 11340 42980
rect 11396 42924 30492 42980
rect 30548 42924 30558 42980
rect 37650 42812 37660 42868
rect 37716 42812 57596 42868
rect 57652 42812 57662 42868
rect 6626 42700 6636 42756
rect 6692 42700 8876 42756
rect 8932 42700 8942 42756
rect 12898 42700 12908 42756
rect 12964 42700 13580 42756
rect 13636 42700 13646 42756
rect 14242 42700 14252 42756
rect 14308 42700 17612 42756
rect 17668 42700 17678 42756
rect 4162 42588 4172 42644
rect 4228 42588 12684 42644
rect 12740 42588 12750 42644
rect 16482 42588 16492 42644
rect 16548 42588 18060 42644
rect 18116 42588 28476 42644
rect 28532 42588 28542 42644
rect 18722 42476 18732 42532
rect 18788 42476 36204 42532
rect 36260 42476 36652 42532
rect 36708 42476 36718 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 7074 42252 7084 42308
rect 7140 42252 11116 42308
rect 11172 42252 11182 42308
rect 23202 42140 23212 42196
rect 23268 42140 24668 42196
rect 24724 42140 27244 42196
rect 27300 42140 27310 42196
rect 29474 42140 29484 42196
rect 29540 42140 31612 42196
rect 31668 42140 31678 42196
rect 31378 42028 31388 42084
rect 31444 42028 33740 42084
rect 33796 42028 33806 42084
rect 40348 42028 45612 42084
rect 45668 42028 45678 42084
rect 40348 41972 40404 42028
rect 14914 41916 14924 41972
rect 14980 41916 16604 41972
rect 16660 41916 16670 41972
rect 37874 41916 37884 41972
rect 37940 41916 40404 41972
rect 41794 41916 41804 41972
rect 41860 41916 44156 41972
rect 44212 41916 44222 41972
rect 41804 41860 41860 41916
rect 728 41832 1820 41860
rect 200 41804 1820 41832
rect 1876 41804 1886 41860
rect 35522 41804 35532 41860
rect 35588 41804 41860 41860
rect 200 41608 800 41804
rect 32610 41692 32620 41748
rect 32676 41692 35420 41748
rect 35476 41692 39676 41748
rect 39732 41692 39742 41748
rect 37538 41580 37548 41636
rect 37604 41580 39900 41636
rect 39956 41580 39966 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 35634 41468 35644 41524
rect 35700 41468 36876 41524
rect 36932 41468 36942 41524
rect 31892 41356 35532 41412
rect 35588 41356 35598 41412
rect 31892 41300 31948 41356
rect 28354 41244 28364 41300
rect 28420 41244 28812 41300
rect 28868 41244 29820 41300
rect 29876 41244 29886 41300
rect 30146 41244 30156 41300
rect 30212 41244 31948 41300
rect 35298 41244 35308 41300
rect 35364 41244 36428 41300
rect 36484 41244 37660 41300
rect 37716 41244 37726 41300
rect 42802 41244 42812 41300
rect 42868 41244 43596 41300
rect 43652 41244 43662 41300
rect 15474 41132 15484 41188
rect 15540 41132 16716 41188
rect 16772 41132 20524 41188
rect 20580 41132 21532 41188
rect 21588 41132 21598 41188
rect 22754 41132 22764 41188
rect 22820 41132 28308 41188
rect 29698 41132 29708 41188
rect 29764 41132 29774 41188
rect 9762 41020 9772 41076
rect 9828 41020 11396 41076
rect 16594 41020 16604 41076
rect 16660 41020 17388 41076
rect 17444 41020 17454 41076
rect 26786 41020 26796 41076
rect 26852 41020 27916 41076
rect 27972 41020 27982 41076
rect 11340 40964 11396 41020
rect 6178 40908 6188 40964
rect 6244 40908 6636 40964
rect 6692 40908 6702 40964
rect 7410 40908 7420 40964
rect 7476 40908 10556 40964
rect 10612 40908 10622 40964
rect 11330 40908 11340 40964
rect 11396 40908 18956 40964
rect 19012 40908 19022 40964
rect 24322 40908 24332 40964
rect 24388 40908 28084 40964
rect 6636 40852 6692 40908
rect 6636 40796 16828 40852
rect 16884 40796 16894 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 28028 40740 28084 40908
rect 28252 40852 28308 41132
rect 29708 41076 29764 41132
rect 59200 41076 59800 41160
rect 29708 41020 29932 41076
rect 29988 41020 35084 41076
rect 35140 41020 35150 41076
rect 35970 41020 35980 41076
rect 36036 41020 38836 41076
rect 39218 41020 39228 41076
rect 39284 41020 43260 41076
rect 43316 41020 43708 41076
rect 57250 41020 57260 41076
rect 57316 41020 58044 41076
rect 58100 41020 59800 41076
rect 38780 40964 38836 41020
rect 43652 40964 43708 41020
rect 31714 40908 31724 40964
rect 31780 40908 33404 40964
rect 33460 40908 33470 40964
rect 34626 40908 34636 40964
rect 34692 40908 37548 40964
rect 37604 40908 38556 40964
rect 38612 40908 38622 40964
rect 38780 40908 40012 40964
rect 40068 40908 40236 40964
rect 40292 40908 40572 40964
rect 40628 40908 40638 40964
rect 43652 40908 43820 40964
rect 43876 40908 48972 40964
rect 49028 40908 49038 40964
rect 59200 40936 59800 41020
rect 28252 40796 37884 40852
rect 37940 40796 37950 40852
rect 38770 40796 38780 40852
rect 38836 40796 40684 40852
rect 40740 40796 42028 40852
rect 42084 40796 42756 40852
rect 42700 40740 42756 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 26338 40684 26348 40740
rect 26404 40684 27804 40740
rect 27860 40684 27870 40740
rect 28028 40684 40460 40740
rect 40516 40684 41132 40740
rect 41188 40684 42140 40740
rect 42196 40684 42206 40740
rect 42690 40684 42700 40740
rect 42756 40684 42766 40740
rect 22194 40572 22204 40628
rect 22260 40572 23660 40628
rect 23716 40572 27692 40628
rect 27748 40572 27758 40628
rect 27906 40572 27916 40628
rect 27972 40572 30044 40628
rect 30100 40572 31052 40628
rect 31108 40572 31118 40628
rect 32050 40572 32060 40628
rect 32116 40572 32620 40628
rect 32676 40572 32686 40628
rect 34850 40572 34860 40628
rect 34916 40572 35980 40628
rect 36036 40572 36046 40628
rect 38546 40572 38556 40628
rect 38612 40572 50876 40628
rect 50932 40572 50942 40628
rect 10546 40460 10556 40516
rect 10612 40460 15148 40516
rect 16594 40460 16604 40516
rect 16660 40460 18620 40516
rect 18676 40460 19068 40516
rect 19124 40460 19628 40516
rect 19684 40460 20636 40516
rect 20692 40460 20702 40516
rect 25890 40460 25900 40516
rect 25956 40460 27244 40516
rect 27300 40460 27468 40516
rect 27524 40460 28476 40516
rect 28532 40460 28542 40516
rect 30482 40460 30492 40516
rect 30548 40460 31164 40516
rect 31220 40460 31230 40516
rect 31826 40460 31836 40516
rect 31892 40460 31902 40516
rect 35074 40460 35084 40516
rect 35140 40460 36204 40516
rect 36260 40460 43372 40516
rect 43428 40460 43438 40516
rect 15092 40404 15148 40460
rect 31836 40404 31892 40460
rect 15092 40348 31892 40404
rect 33842 40348 33852 40404
rect 33908 40348 34972 40404
rect 35028 40348 35980 40404
rect 36036 40348 36046 40404
rect 36530 40348 36540 40404
rect 36596 40348 38780 40404
rect 38836 40348 38846 40404
rect 40226 40348 40236 40404
rect 40292 40348 41468 40404
rect 41524 40348 57708 40404
rect 57764 40348 57774 40404
rect 19730 40236 19740 40292
rect 19796 40236 23212 40292
rect 23268 40236 23278 40292
rect 26898 40236 26908 40292
rect 26964 40236 27356 40292
rect 27412 40236 28140 40292
rect 28196 40236 28364 40292
rect 28420 40236 28430 40292
rect 29698 40236 29708 40292
rect 29764 40236 31836 40292
rect 31892 40236 31902 40292
rect 33058 40236 33068 40292
rect 33124 40236 34300 40292
rect 34356 40236 36652 40292
rect 36708 40236 36718 40292
rect 42466 40236 42476 40292
rect 42532 40236 43148 40292
rect 43204 40236 43214 40292
rect 47618 40236 47628 40292
rect 47684 40236 48188 40292
rect 48244 40236 48254 40292
rect 20738 40124 20748 40180
rect 20804 40124 24220 40180
rect 24276 40124 33908 40180
rect 34066 40124 34076 40180
rect 34132 40124 34748 40180
rect 34804 40124 34814 40180
rect 34972 40124 40796 40180
rect 40852 40124 40862 40180
rect 33852 40068 33908 40124
rect 34972 40068 35028 40124
rect 42476 40068 42532 40236
rect 24098 40012 24108 40068
rect 24164 40012 33180 40068
rect 33236 40012 33246 40068
rect 33852 40012 35028 40068
rect 35634 40012 35644 40068
rect 35700 40012 37548 40068
rect 37604 40012 40684 40068
rect 40740 40012 42532 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 7186 39900 7196 39956
rect 7252 39900 34524 39956
rect 34580 39900 34590 39956
rect 20066 39788 20076 39844
rect 20132 39788 34636 39844
rect 34692 39788 34702 39844
rect 38546 39788 38556 39844
rect 38612 39788 40572 39844
rect 40628 39788 41804 39844
rect 41860 39788 41870 39844
rect 36418 39676 36428 39732
rect 36484 39676 38332 39732
rect 38388 39676 38398 39732
rect 19506 39564 19516 39620
rect 19572 39564 21532 39620
rect 21588 39564 27356 39620
rect 27412 39564 27422 39620
rect 35074 39564 35084 39620
rect 35140 39564 38108 39620
rect 38164 39564 38174 39620
rect 39890 39564 39900 39620
rect 39956 39564 40572 39620
rect 40628 39564 40638 39620
rect 42802 39564 42812 39620
rect 42868 39564 47516 39620
rect 47572 39564 47582 39620
rect 3938 39452 3948 39508
rect 4004 39452 17164 39508
rect 17220 39452 17230 39508
rect 31266 39452 31276 39508
rect 31332 39452 32284 39508
rect 32340 39452 38780 39508
rect 38836 39452 39228 39508
rect 39284 39452 39294 39508
rect 46722 39452 46732 39508
rect 46788 39452 47292 39508
rect 47348 39452 47628 39508
rect 47684 39452 47694 39508
rect 47842 39452 47852 39508
rect 47908 39452 48748 39508
rect 48804 39452 49644 39508
rect 49700 39452 49710 39508
rect 26002 39340 26012 39396
rect 26068 39340 26348 39396
rect 26404 39340 26796 39396
rect 26852 39340 26862 39396
rect 34514 39340 34524 39396
rect 34580 39340 35084 39396
rect 35140 39340 35756 39396
rect 35812 39340 36540 39396
rect 36596 39340 36606 39396
rect 40674 39340 40684 39396
rect 40740 39340 41580 39396
rect 41636 39340 45500 39396
rect 45556 39340 45566 39396
rect 33170 39228 33180 39284
rect 33236 39228 33740 39284
rect 33796 39228 35644 39284
rect 35700 39228 35710 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 23762 39116 23772 39172
rect 23828 39116 35756 39172
rect 35812 39116 36204 39172
rect 36260 39116 36270 39172
rect 4806 39004 4844 39060
rect 4900 39004 4910 39060
rect 17042 39004 17052 39060
rect 17108 39004 20412 39060
rect 20468 39004 21756 39060
rect 21812 39004 21822 39060
rect 27010 39004 27020 39060
rect 27076 39004 27580 39060
rect 27636 39004 27646 39060
rect 30146 39004 30156 39060
rect 30212 39004 30940 39060
rect 30996 39004 31006 39060
rect 45490 39004 45500 39060
rect 45556 39004 46620 39060
rect 46676 39004 46686 39060
rect 12674 38892 12684 38948
rect 12740 38892 13244 38948
rect 13300 38892 31948 38948
rect 32004 38892 32014 38948
rect 36306 38892 36316 38948
rect 36372 38892 39116 38948
rect 39172 38892 39182 38948
rect 40562 38892 40572 38948
rect 40628 38892 41916 38948
rect 41972 38892 41982 38948
rect 23202 38780 23212 38836
rect 23268 38780 45388 38836
rect 45444 38780 45454 38836
rect 45938 38780 45948 38836
rect 46004 38780 48524 38836
rect 48580 38780 48590 38836
rect 3826 38668 3836 38724
rect 3892 38668 4396 38724
rect 4452 38668 4462 38724
rect 36082 38668 36092 38724
rect 36148 38668 38556 38724
rect 38612 38668 38622 38724
rect 40898 38668 40908 38724
rect 40964 38668 41580 38724
rect 41636 38668 41646 38724
rect 43698 38668 43708 38724
rect 43764 38668 44604 38724
rect 44660 38668 45724 38724
rect 45780 38668 45790 38724
rect 3938 38556 3948 38612
rect 4004 38556 8204 38612
rect 8260 38556 8270 38612
rect 35858 38556 35868 38612
rect 35924 38556 36652 38612
rect 36708 38556 36718 38612
rect 200 38276 800 38472
rect 5058 38444 5068 38500
rect 5124 38444 10892 38500
rect 10948 38444 10958 38500
rect 26450 38444 26460 38500
rect 26516 38444 26908 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 26852 38388 26908 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 4834 38332 4844 38388
rect 4900 38332 11340 38388
rect 11396 38332 11406 38388
rect 26852 38332 27804 38388
rect 27860 38332 28812 38388
rect 28868 38332 34468 38388
rect 200 38248 1820 38276
rect 728 38220 1820 38248
rect 1876 38220 1886 38276
rect 12002 38220 12012 38276
rect 12068 38220 16492 38276
rect 16548 38220 16558 38276
rect 27346 38220 27356 38276
rect 27412 38220 30492 38276
rect 30548 38220 30558 38276
rect 34412 38164 34468 38332
rect 13682 38108 13692 38164
rect 13748 38108 14028 38164
rect 14084 38108 24556 38164
rect 24612 38108 25676 38164
rect 25732 38108 32508 38164
rect 32564 38108 32574 38164
rect 34402 38108 34412 38164
rect 34468 38108 35084 38164
rect 35140 38108 35150 38164
rect 41122 38108 41132 38164
rect 41188 38108 41692 38164
rect 41748 38108 41758 38164
rect 12786 37996 12796 38052
rect 12852 37996 13356 38052
rect 13412 37996 13422 38052
rect 17266 37996 17276 38052
rect 17332 37996 18172 38052
rect 18228 37996 18238 38052
rect 24098 37996 24108 38052
rect 24164 37996 25564 38052
rect 25620 37996 25630 38052
rect 26114 37996 26124 38052
rect 26180 37996 26684 38052
rect 26740 37996 26750 38052
rect 31490 37996 31500 38052
rect 31556 37996 32844 38052
rect 32900 37996 32910 38052
rect 33954 37996 33964 38052
rect 34020 37996 35308 38052
rect 35364 37996 35374 38052
rect 39778 37996 39788 38052
rect 39844 37996 42140 38052
rect 42196 37996 43708 38052
rect 43652 37940 43708 37996
rect 12898 37884 12908 37940
rect 12964 37884 13692 37940
rect 13748 37884 13758 37940
rect 14242 37884 14252 37940
rect 14308 37884 25900 37940
rect 25956 37884 27356 37940
rect 27412 37884 27422 37940
rect 30370 37884 30380 37940
rect 30436 37884 31948 37940
rect 32004 37884 32014 37940
rect 38434 37884 38444 37940
rect 38500 37884 39116 37940
rect 39172 37884 39182 37940
rect 43652 37884 57596 37940
rect 57652 37884 57662 37940
rect 14578 37772 14588 37828
rect 14644 37772 15596 37828
rect 15652 37772 23100 37828
rect 23156 37772 25004 37828
rect 25060 37772 26124 37828
rect 26180 37772 26190 37828
rect 39414 37772 39452 37828
rect 39508 37772 39518 37828
rect 57250 37772 57260 37828
rect 57316 37772 58044 37828
rect 58100 37800 59304 37828
rect 58100 37772 59800 37800
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37576 59800 37772
rect 16930 37436 16940 37492
rect 16996 37436 17724 37492
rect 17780 37436 17790 37492
rect 18946 37436 18956 37492
rect 19012 37436 19068 37492
rect 19124 37436 19134 37492
rect 19282 37436 19292 37492
rect 19348 37436 20524 37492
rect 20580 37436 32060 37492
rect 32116 37436 32126 37492
rect 32582 37436 32620 37492
rect 32676 37436 33180 37492
rect 33236 37436 33246 37492
rect 36194 37436 36204 37492
rect 36260 37436 36652 37492
rect 36708 37436 36718 37492
rect 42466 37436 42476 37492
rect 42532 37436 43484 37492
rect 43540 37436 57708 37492
rect 57764 37436 57774 37492
rect 11778 37324 11788 37380
rect 11844 37324 13132 37380
rect 13188 37324 24108 37380
rect 24164 37324 24174 37380
rect 24994 37324 25004 37380
rect 25060 37324 25788 37380
rect 25844 37324 25854 37380
rect 26236 37324 27244 37380
rect 27300 37324 27310 37380
rect 30930 37324 30940 37380
rect 30996 37324 31276 37380
rect 31332 37324 31500 37380
rect 31556 37324 31566 37380
rect 10882 37212 10892 37268
rect 10948 37212 12572 37268
rect 12628 37212 12638 37268
rect 18834 37212 18844 37268
rect 18900 37212 19180 37268
rect 19236 37212 19246 37268
rect 19730 37212 19740 37268
rect 19796 37212 20972 37268
rect 21028 37212 25676 37268
rect 25732 37212 25742 37268
rect 26236 37156 26292 37324
rect 26898 37212 26908 37268
rect 26964 37212 28812 37268
rect 28868 37212 33964 37268
rect 34020 37212 34030 37268
rect 40450 37212 40460 37268
rect 40516 37212 41468 37268
rect 41524 37212 41534 37268
rect 11442 37100 11452 37156
rect 11508 37100 13020 37156
rect 13076 37100 13086 37156
rect 13234 37100 13244 37156
rect 13300 37100 15036 37156
rect 15092 37100 15372 37156
rect 15428 37100 26292 37156
rect 31938 37100 31948 37156
rect 32004 37100 35084 37156
rect 35140 37100 41132 37156
rect 41188 37100 41198 37156
rect 18498 36988 18508 37044
rect 18564 36988 18732 37044
rect 18788 36988 19964 37044
rect 20020 36988 20030 37044
rect 25666 36988 25676 37044
rect 25732 36988 26572 37044
rect 26628 36988 29148 37044
rect 29204 36988 29214 37044
rect 33170 36988 33180 37044
rect 33236 36988 35868 37044
rect 35924 36988 35934 37044
rect 48636 36988 49980 37044
rect 50036 36988 50988 37044
rect 51044 36988 51054 37044
rect 48636 36932 48692 36988
rect 12002 36876 12012 36932
rect 12068 36876 12684 36932
rect 12740 36876 12750 36932
rect 13458 36876 13468 36932
rect 13524 36876 14028 36932
rect 14084 36876 14094 36932
rect 17154 36876 17164 36932
rect 17220 36876 17724 36932
rect 17780 36876 17790 36932
rect 23538 36876 23548 36932
rect 23604 36876 24444 36932
rect 24500 36876 24510 36932
rect 39778 36876 39788 36932
rect 39844 36876 41692 36932
rect 41748 36876 41758 36932
rect 41906 36876 41916 36932
rect 41972 36876 46060 36932
rect 46116 36876 48692 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 7970 36764 7980 36820
rect 8036 36764 32284 36820
rect 32340 36764 32732 36820
rect 32788 36764 32798 36820
rect 35634 36764 35644 36820
rect 35700 36764 43036 36820
rect 43092 36764 43102 36820
rect 3602 36652 3612 36708
rect 3668 36652 3836 36708
rect 3892 36652 5628 36708
rect 5684 36652 5694 36708
rect 8978 36652 8988 36708
rect 9044 36652 11900 36708
rect 11956 36652 11966 36708
rect 12450 36652 12460 36708
rect 12516 36652 13244 36708
rect 13300 36652 13310 36708
rect 17938 36652 17948 36708
rect 18004 36652 32732 36708
rect 32788 36652 32798 36708
rect 33506 36652 33516 36708
rect 33572 36652 34076 36708
rect 34132 36652 34972 36708
rect 35028 36652 35038 36708
rect 40562 36652 40572 36708
rect 40628 36652 41356 36708
rect 41412 36652 41422 36708
rect 4050 36540 4060 36596
rect 4116 36540 8876 36596
rect 8932 36540 8942 36596
rect 17350 36540 17388 36596
rect 17444 36540 17454 36596
rect 19030 36540 19068 36596
rect 19124 36540 19134 36596
rect 19842 36540 19852 36596
rect 19908 36540 20412 36596
rect 20468 36540 32452 36596
rect 34402 36540 34412 36596
rect 34468 36540 34860 36596
rect 34916 36540 35532 36596
rect 35588 36540 36540 36596
rect 36596 36540 37212 36596
rect 37268 36540 37278 36596
rect 41570 36540 41580 36596
rect 41636 36540 42140 36596
rect 42196 36540 42206 36596
rect 32396 36484 32452 36540
rect 3490 36428 3500 36484
rect 3556 36428 6412 36484
rect 6468 36428 7308 36484
rect 7364 36428 7374 36484
rect 11442 36428 11452 36484
rect 11508 36428 11900 36484
rect 11956 36428 11966 36484
rect 14130 36428 14140 36484
rect 14196 36428 15148 36484
rect 15204 36428 15214 36484
rect 17826 36428 17836 36484
rect 17892 36428 19180 36484
rect 19236 36428 19246 36484
rect 19394 36428 19404 36484
rect 19460 36428 25116 36484
rect 25172 36428 25182 36484
rect 30594 36428 30604 36484
rect 30660 36428 31388 36484
rect 31444 36428 32172 36484
rect 32228 36428 32238 36484
rect 32396 36428 33012 36484
rect 33506 36428 33516 36484
rect 33572 36428 34076 36484
rect 34132 36428 34636 36484
rect 34692 36428 34702 36484
rect 35970 36428 35980 36484
rect 36036 36428 40124 36484
rect 40180 36428 40190 36484
rect 41122 36428 41132 36484
rect 41188 36428 43708 36484
rect 43764 36428 45164 36484
rect 45220 36428 45230 36484
rect 19404 36372 19460 36428
rect 32956 36372 33012 36428
rect 41132 36372 41188 36428
rect 4386 36316 4396 36372
rect 4452 36316 5068 36372
rect 5124 36316 7532 36372
rect 7588 36316 8652 36372
rect 8708 36316 8718 36372
rect 12786 36316 12796 36372
rect 12852 36316 13468 36372
rect 13524 36316 13534 36372
rect 16482 36316 16492 36372
rect 16548 36316 18284 36372
rect 18340 36316 19460 36372
rect 24098 36316 24108 36372
rect 24164 36316 24892 36372
rect 24948 36316 25228 36372
rect 25284 36316 25294 36372
rect 32956 36316 37100 36372
rect 37156 36316 37166 36372
rect 37426 36316 37436 36372
rect 37492 36316 40012 36372
rect 40068 36316 41188 36372
rect 4498 36204 4508 36260
rect 4564 36204 8764 36260
rect 8820 36204 8830 36260
rect 9202 36204 9212 36260
rect 9268 36204 10108 36260
rect 10164 36204 11900 36260
rect 11956 36204 11966 36260
rect 16034 36204 16044 36260
rect 16100 36204 16716 36260
rect 16772 36204 16782 36260
rect 17826 36204 17836 36260
rect 17892 36204 18060 36260
rect 18116 36204 18732 36260
rect 18788 36204 18956 36260
rect 19012 36204 20188 36260
rect 20244 36204 20254 36260
rect 22866 36204 22876 36260
rect 22932 36204 23548 36260
rect 23604 36204 23614 36260
rect 24770 36204 24780 36260
rect 24836 36204 26572 36260
rect 26628 36204 29708 36260
rect 29764 36204 30044 36260
rect 30100 36204 30380 36260
rect 30436 36204 30446 36260
rect 32834 36204 32844 36260
rect 32900 36204 38668 36260
rect 39554 36204 39564 36260
rect 39620 36204 40684 36260
rect 40740 36204 40750 36260
rect 38612 36148 38668 36204
rect 19142 36092 19180 36148
rect 19236 36092 19246 36148
rect 26852 36092 35644 36148
rect 35700 36092 35710 36148
rect 38612 36092 39676 36148
rect 39732 36092 39742 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26852 36036 26908 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4722 35980 4732 36036
rect 4788 35980 5292 36036
rect 5348 35980 9884 36036
rect 9940 35980 9950 36036
rect 12012 35980 12236 36036
rect 12292 35980 12302 36036
rect 14466 35980 14476 36036
rect 14532 35980 16044 36036
rect 16100 35980 16110 36036
rect 25666 35980 25676 36036
rect 25732 35980 26236 36036
rect 26292 35980 26908 36036
rect 33618 35980 33628 36036
rect 33684 35980 34860 36036
rect 34916 35980 35980 36036
rect 36036 35980 36046 36036
rect 12012 35924 12068 35980
rect 3378 35868 3388 35924
rect 3444 35868 8204 35924
rect 8260 35868 10108 35924
rect 10164 35868 10174 35924
rect 12002 35868 12012 35924
rect 12068 35868 12078 35924
rect 12562 35868 12572 35924
rect 12628 35868 14140 35924
rect 14196 35868 14206 35924
rect 14354 35868 14364 35924
rect 14420 35868 14700 35924
rect 14756 35868 17500 35924
rect 17556 35868 17566 35924
rect 19282 35868 19292 35924
rect 19348 35868 20076 35924
rect 20132 35868 20142 35924
rect 21746 35868 21756 35924
rect 21812 35868 45948 35924
rect 46004 35868 46014 35924
rect 728 35784 1708 35812
rect 200 35756 1708 35784
rect 1764 35756 1774 35812
rect 6850 35756 6860 35812
rect 6916 35756 7980 35812
rect 8036 35756 9212 35812
rect 9268 35756 9772 35812
rect 9828 35756 9838 35812
rect 12236 35756 12460 35812
rect 12516 35756 12908 35812
rect 12964 35756 15372 35812
rect 15428 35756 16492 35812
rect 16548 35756 16558 35812
rect 18274 35756 18284 35812
rect 18340 35756 19852 35812
rect 19908 35756 29708 35812
rect 29764 35756 29932 35812
rect 29988 35756 30716 35812
rect 30772 35756 30782 35812
rect 33170 35756 33180 35812
rect 33236 35756 33628 35812
rect 33684 35756 33694 35812
rect 34962 35756 34972 35812
rect 35028 35756 35644 35812
rect 35700 35756 35710 35812
rect 37090 35756 37100 35812
rect 37156 35756 38220 35812
rect 38276 35756 39564 35812
rect 39620 35756 39630 35812
rect 44706 35756 44716 35812
rect 44772 35756 45836 35812
rect 45892 35756 45902 35812
rect 46050 35756 46060 35812
rect 46116 35756 47292 35812
rect 47348 35756 47358 35812
rect 200 35560 800 35756
rect 12236 35700 12292 35756
rect 12226 35644 12236 35700
rect 12292 35644 12302 35700
rect 15474 35644 15484 35700
rect 15540 35644 16268 35700
rect 16324 35644 16828 35700
rect 16884 35644 16894 35700
rect 17826 35644 17836 35700
rect 17892 35644 19292 35700
rect 19348 35644 19358 35700
rect 32386 35644 32396 35700
rect 32452 35644 34188 35700
rect 34244 35644 34412 35700
rect 34468 35644 34478 35700
rect 45154 35644 45164 35700
rect 45220 35644 46284 35700
rect 46340 35644 46350 35700
rect 46498 35644 46508 35700
rect 46564 35644 49420 35700
rect 49476 35644 49486 35700
rect 50082 35644 50092 35700
rect 50148 35644 50876 35700
rect 50932 35644 51884 35700
rect 51940 35644 51950 35700
rect 6300 35532 13356 35588
rect 13412 35532 14028 35588
rect 14084 35532 14094 35588
rect 15138 35532 15148 35588
rect 15204 35532 26012 35588
rect 26068 35532 26078 35588
rect 32834 35532 32844 35588
rect 32900 35532 33740 35588
rect 33796 35532 33806 35588
rect 35746 35532 35756 35588
rect 35812 35532 36652 35588
rect 36708 35532 38668 35588
rect 38724 35532 39788 35588
rect 39844 35532 39854 35588
rect 40002 35532 40012 35588
rect 40068 35532 40078 35588
rect 6300 35476 6356 35532
rect 3490 35420 3500 35476
rect 3556 35420 6300 35476
rect 6356 35420 6366 35476
rect 10434 35420 10444 35476
rect 10500 35420 11340 35476
rect 11396 35420 11676 35476
rect 11732 35420 16716 35476
rect 16772 35420 24892 35476
rect 24948 35420 24958 35476
rect 31490 35420 31500 35476
rect 31556 35420 38108 35476
rect 38164 35420 38174 35476
rect 5506 35308 5516 35364
rect 5572 35308 8988 35364
rect 9044 35308 9548 35364
rect 9604 35308 9614 35364
rect 16034 35308 16044 35364
rect 16100 35308 16940 35364
rect 16996 35308 17836 35364
rect 17892 35308 18060 35364
rect 18116 35308 18126 35364
rect 18274 35308 18284 35364
rect 18340 35308 18350 35364
rect 19506 35308 19516 35364
rect 19572 35308 19582 35364
rect 25442 35308 25452 35364
rect 25508 35308 26236 35364
rect 26292 35308 26302 35364
rect 35858 35308 35868 35364
rect 35924 35308 36316 35364
rect 36372 35308 36652 35364
rect 36708 35308 36718 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 18284 35252 18340 35308
rect 12562 35196 12572 35252
rect 12628 35196 15820 35252
rect 15876 35196 15886 35252
rect 17266 35196 17276 35252
rect 17332 35196 18340 35252
rect 19516 35252 19572 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 40012 35252 40068 35532
rect 43652 35420 51324 35476
rect 51380 35420 51390 35476
rect 43652 35364 43708 35420
rect 41794 35308 41804 35364
rect 41860 35308 43708 35364
rect 19516 35196 22540 35252
rect 22596 35196 22606 35252
rect 22764 35196 29148 35252
rect 29204 35196 29214 35252
rect 29362 35196 29372 35252
rect 29428 35196 30156 35252
rect 30212 35196 34972 35252
rect 35028 35196 35038 35252
rect 39106 35196 39116 35252
rect 39172 35196 40068 35252
rect 40562 35196 40572 35252
rect 40628 35196 49308 35252
rect 49364 35196 49532 35252
rect 49588 35196 49980 35252
rect 50036 35196 50046 35252
rect 22764 35140 22820 35196
rect 8530 35084 8540 35140
rect 8596 35084 11340 35140
rect 11396 35084 11564 35140
rect 11620 35084 11630 35140
rect 22092 35084 22820 35140
rect 24994 35084 25004 35140
rect 25060 35084 26908 35140
rect 26964 35084 29596 35140
rect 29652 35084 29662 35140
rect 36306 35084 36316 35140
rect 36372 35084 40236 35140
rect 40292 35084 40302 35140
rect 22092 34916 22148 35084
rect 59200 35028 59800 35112
rect 22418 34972 22428 35028
rect 22484 34972 22988 35028
rect 23044 34972 39452 35028
rect 39508 34972 39518 35028
rect 42690 34972 42700 35028
rect 42756 34972 43148 35028
rect 43204 34972 44716 35028
rect 44772 34972 45164 35028
rect 45220 34972 45230 35028
rect 52882 34972 52892 35028
rect 52948 34972 56252 35028
rect 56308 34972 56812 35028
rect 56868 34972 56878 35028
rect 57810 34972 57820 35028
rect 57876 34972 59800 35028
rect 20402 34860 20412 34916
rect 20468 34860 22092 34916
rect 22148 34860 22158 34916
rect 24994 34860 25004 34916
rect 25060 34860 26348 34916
rect 26404 34860 26414 34916
rect 29138 34860 29148 34916
rect 29204 34860 36876 34916
rect 36932 34860 36942 34916
rect 59200 34888 59800 34972
rect 9090 34748 9100 34804
rect 9156 34748 10220 34804
rect 10276 34748 10286 34804
rect 10770 34748 10780 34804
rect 10836 34748 11788 34804
rect 11844 34748 12572 34804
rect 12628 34748 12638 34804
rect 18498 34748 18508 34804
rect 18564 34748 19068 34804
rect 19124 34748 19134 34804
rect 25442 34748 25452 34804
rect 25508 34748 26684 34804
rect 26740 34748 26750 34804
rect 9986 34636 9996 34692
rect 10052 34636 10332 34692
rect 10388 34636 10398 34692
rect 15810 34636 15820 34692
rect 15876 34636 19292 34692
rect 19348 34636 19852 34692
rect 19908 34636 20244 34692
rect 20850 34636 20860 34692
rect 20916 34636 21980 34692
rect 22036 34636 22046 34692
rect 24210 34636 24220 34692
rect 24276 34636 25228 34692
rect 25284 34636 25294 34692
rect 35074 34636 35084 34692
rect 35140 34636 36092 34692
rect 36148 34636 36158 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 20188 34468 20244 34636
rect 21746 34524 21756 34580
rect 21812 34524 23324 34580
rect 23380 34524 29484 34580
rect 29540 34524 29550 34580
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 20188 34412 27916 34468
rect 27972 34412 27982 34468
rect 28466 34412 28476 34468
rect 28532 34412 36988 34468
rect 37044 34412 39116 34468
rect 39172 34412 39182 34468
rect 45938 34412 45948 34468
rect 46004 34412 46732 34468
rect 46788 34412 46798 34468
rect 7970 34300 7980 34356
rect 8036 34300 8540 34356
rect 8596 34300 8606 34356
rect 10546 34300 10556 34356
rect 10612 34300 11228 34356
rect 11284 34300 11294 34356
rect 34962 34300 34972 34356
rect 35028 34300 35868 34356
rect 35924 34300 36092 34356
rect 36148 34300 36158 34356
rect 45154 34300 45164 34356
rect 45220 34300 45836 34356
rect 45892 34300 45902 34356
rect 2146 34188 2156 34244
rect 2212 34188 4732 34244
rect 4788 34188 4798 34244
rect 8082 34188 8092 34244
rect 8148 34188 8876 34244
rect 8932 34188 10444 34244
rect 10500 34188 10510 34244
rect 20514 34188 20524 34244
rect 20580 34188 23772 34244
rect 23828 34188 25676 34244
rect 25732 34188 25742 34244
rect 26338 34188 26348 34244
rect 26404 34188 39900 34244
rect 39956 34188 39966 34244
rect 9874 34076 9884 34132
rect 9940 34076 10668 34132
rect 10724 34076 11228 34132
rect 11284 34076 11294 34132
rect 23874 34076 23884 34132
rect 23940 34076 25116 34132
rect 25172 34076 29708 34132
rect 29764 34076 29774 34132
rect 33842 34076 33852 34132
rect 33908 34076 34636 34132
rect 34692 34076 34702 34132
rect 38612 34076 40572 34132
rect 40628 34076 40638 34132
rect 38612 34020 38668 34076
rect 4946 33964 4956 34020
rect 5012 33964 9772 34020
rect 9828 33964 9838 34020
rect 19394 33964 19404 34020
rect 19460 33964 19852 34020
rect 19908 33964 20412 34020
rect 20468 33964 20478 34020
rect 26114 33964 26124 34020
rect 26180 33964 26572 34020
rect 26628 33964 26638 34020
rect 27906 33964 27916 34020
rect 27972 33964 36764 34020
rect 36820 33964 36988 34020
rect 37044 33964 38668 34020
rect 26572 33908 26628 33964
rect 8642 33852 8652 33908
rect 8708 33852 10220 33908
rect 10276 33852 11676 33908
rect 11732 33852 15148 33908
rect 19954 33852 19964 33908
rect 20020 33852 20188 33908
rect 20244 33852 21644 33908
rect 21700 33852 21710 33908
rect 26572 33852 39228 33908
rect 39284 33852 39294 33908
rect 9426 33740 9436 33796
rect 9492 33740 9996 33796
rect 10052 33740 10062 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 15092 33684 15148 33852
rect 26852 33740 28476 33796
rect 28532 33740 28542 33796
rect 15092 33628 20300 33684
rect 20356 33628 20366 33684
rect 25218 33628 25228 33684
rect 25284 33628 26796 33684
rect 26852 33628 26908 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 10770 33516 10780 33572
rect 10836 33516 11452 33572
rect 11508 33516 34076 33572
rect 34132 33516 34142 33572
rect 34850 33516 34860 33572
rect 34916 33516 38332 33572
rect 38388 33516 38398 33572
rect 11218 33404 11228 33460
rect 11284 33404 11900 33460
rect 11956 33404 11966 33460
rect 17154 33404 17164 33460
rect 17220 33404 17612 33460
rect 17668 33404 17678 33460
rect 23986 33404 23996 33460
rect 24052 33404 25452 33460
rect 25508 33404 26012 33460
rect 26068 33404 26078 33460
rect 29698 33404 29708 33460
rect 29764 33404 30268 33460
rect 30324 33404 30334 33460
rect 36418 33404 36428 33460
rect 36484 33404 42028 33460
rect 42084 33404 42476 33460
rect 42532 33404 42542 33460
rect 8642 33292 8652 33348
rect 8708 33292 18844 33348
rect 18900 33292 18910 33348
rect 22306 33292 22316 33348
rect 22372 33292 24444 33348
rect 24500 33292 25788 33348
rect 25844 33292 25854 33348
rect 35410 33292 35420 33348
rect 35476 33292 35644 33348
rect 35700 33292 40908 33348
rect 40964 33292 41916 33348
rect 41972 33292 41982 33348
rect 11890 33180 11900 33236
rect 11956 33180 18620 33236
rect 18676 33180 18686 33236
rect 27794 33180 27804 33236
rect 27860 33180 28028 33236
rect 28084 33180 28252 33236
rect 28308 33180 28318 33236
rect 28914 33180 28924 33236
rect 28980 33180 29596 33236
rect 29652 33180 29662 33236
rect 36642 33180 36652 33236
rect 36708 33180 37324 33236
rect 37380 33180 38892 33236
rect 38948 33180 38958 33236
rect 19282 33068 19292 33124
rect 19348 33068 25004 33124
rect 25060 33068 25564 33124
rect 25620 33068 25630 33124
rect 27468 33068 27692 33124
rect 27748 33068 27758 33124
rect 35522 33068 35532 33124
rect 35588 33068 36092 33124
rect 36148 33068 36158 33124
rect 41682 33068 41692 33124
rect 41748 33068 50092 33124
rect 50148 33068 50316 33124
rect 50372 33068 50540 33124
rect 50596 33068 57708 33124
rect 57764 33068 57774 33124
rect 27468 33012 27524 33068
rect 9650 32956 9660 33012
rect 9716 32956 10164 33012
rect 26758 32956 26796 33012
rect 26852 32956 26862 33012
rect 27458 32956 27468 33012
rect 27524 32956 27534 33012
rect 29474 32956 29484 33012
rect 29540 32956 32508 33012
rect 32564 32956 33068 33012
rect 33124 32956 38220 33012
rect 38276 32956 39004 33012
rect 39060 32956 39070 33012
rect 10108 32788 10164 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 27234 32844 27244 32900
rect 27300 32844 28588 32900
rect 28644 32844 37100 32900
rect 37156 32844 37166 32900
rect 10108 32732 11452 32788
rect 11508 32732 11518 32788
rect 26898 32732 26908 32788
rect 26964 32732 27636 32788
rect 33954 32732 33964 32788
rect 34020 32732 34524 32788
rect 34580 32732 34590 32788
rect 35186 32732 35196 32788
rect 35252 32732 37212 32788
rect 37268 32732 37884 32788
rect 37940 32732 37950 32788
rect 10108 32564 10164 32732
rect 27580 32676 27636 32732
rect 10882 32620 10892 32676
rect 10948 32620 11564 32676
rect 11620 32620 12292 32676
rect 12450 32620 12460 32676
rect 12516 32620 13580 32676
rect 13636 32620 15148 32676
rect 15204 32620 15214 32676
rect 25666 32620 25676 32676
rect 25732 32620 27244 32676
rect 27300 32620 27310 32676
rect 27570 32620 27580 32676
rect 27636 32620 27646 32676
rect 39890 32620 39900 32676
rect 39956 32620 42700 32676
rect 42756 32620 42766 32676
rect 12236 32564 12292 32620
rect 10098 32508 10108 32564
rect 10164 32508 10174 32564
rect 12226 32508 12236 32564
rect 12292 32508 12302 32564
rect 21410 32508 21420 32564
rect 21476 32508 22204 32564
rect 22260 32508 22270 32564
rect 24994 32508 25004 32564
rect 25060 32508 26236 32564
rect 26292 32508 28924 32564
rect 28980 32508 28990 32564
rect 728 32424 2044 32452
rect 200 32396 2044 32424
rect 2100 32396 2110 32452
rect 12562 32396 12572 32452
rect 12628 32396 13132 32452
rect 13188 32396 13198 32452
rect 22642 32396 22652 32452
rect 22708 32396 23772 32452
rect 23828 32396 32060 32452
rect 32116 32396 35196 32452
rect 35252 32396 35868 32452
rect 35924 32396 35934 32452
rect 36978 32396 36988 32452
rect 37044 32396 40124 32452
rect 40180 32396 40190 32452
rect 200 32200 800 32396
rect 22866 32284 22876 32340
rect 22932 32284 23324 32340
rect 23380 32284 24108 32340
rect 24164 32284 26012 32340
rect 26068 32284 29372 32340
rect 29428 32284 29438 32340
rect 38434 32284 38444 32340
rect 38500 32284 40684 32340
rect 40740 32284 40750 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 27244 32116 27300 32284
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 7858 32060 7868 32116
rect 7924 32060 9772 32116
rect 9828 32060 11004 32116
rect 11060 32060 11070 32116
rect 27234 32060 27244 32116
rect 27300 32060 27310 32116
rect 38994 32060 39004 32116
rect 39060 32060 39900 32116
rect 39956 32060 39966 32116
rect 13010 31948 13020 32004
rect 13076 31948 13916 32004
rect 13972 31948 13982 32004
rect 40002 31948 40012 32004
rect 40068 31948 40348 32004
rect 40404 31948 40414 32004
rect 5618 31836 5628 31892
rect 5684 31836 6412 31892
rect 6468 31836 6478 31892
rect 10434 31836 10444 31892
rect 10500 31836 11004 31892
rect 11060 31836 11070 31892
rect 11890 31836 11900 31892
rect 11956 31836 12124 31892
rect 12180 31836 12190 31892
rect 16034 31836 16044 31892
rect 16100 31836 17052 31892
rect 17108 31836 17118 31892
rect 28130 31836 28140 31892
rect 28196 31836 30492 31892
rect 30548 31836 30558 31892
rect 38658 31836 38668 31892
rect 38724 31836 39228 31892
rect 39284 31836 39294 31892
rect 11676 31724 11788 31780
rect 11844 31724 11854 31780
rect 20962 31724 20972 31780
rect 21028 31724 26908 31780
rect 29922 31724 29932 31780
rect 29988 31724 36876 31780
rect 36932 31724 38108 31780
rect 38164 31724 38174 31780
rect 11676 31556 11732 31724
rect 26852 31668 26908 31724
rect 11890 31612 11900 31668
rect 11956 31612 12684 31668
rect 12740 31612 12750 31668
rect 13906 31612 13916 31668
rect 13972 31612 16604 31668
rect 16660 31612 18060 31668
rect 18116 31612 18126 31668
rect 26852 31612 37772 31668
rect 37828 31612 37838 31668
rect 39442 31612 39452 31668
rect 39508 31612 40348 31668
rect 40404 31612 40414 31668
rect 59200 31556 59800 31752
rect 11666 31500 11676 31556
rect 11732 31500 12348 31556
rect 12404 31500 12414 31556
rect 23874 31500 23884 31556
rect 23940 31500 24332 31556
rect 24388 31500 24398 31556
rect 37874 31500 37884 31556
rect 37940 31500 39564 31556
rect 39620 31500 40460 31556
rect 40516 31500 41356 31556
rect 41412 31500 42140 31556
rect 42196 31500 42206 31556
rect 58034 31500 58044 31556
rect 58100 31528 59800 31556
rect 58100 31500 59304 31528
rect 6402 31388 6412 31444
rect 6468 31388 16044 31444
rect 16100 31388 16380 31444
rect 16436 31388 16446 31444
rect 26852 31388 30604 31444
rect 30660 31388 31724 31444
rect 31780 31388 36204 31444
rect 36260 31388 39900 31444
rect 39956 31388 40124 31444
rect 40180 31388 40572 31444
rect 40628 31388 40638 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 8530 31276 8540 31332
rect 8596 31276 15148 31332
rect 15092 31220 15148 31276
rect 26852 31220 26908 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 10882 31164 10892 31220
rect 10948 31164 11340 31220
rect 11396 31164 12068 31220
rect 15092 31164 23660 31220
rect 23716 31164 24780 31220
rect 24836 31164 26908 31220
rect 30818 31164 30828 31220
rect 30884 31164 31276 31220
rect 31332 31164 57484 31220
rect 57540 31164 57550 31220
rect 12012 31108 12068 31164
rect 12002 31052 12012 31108
rect 12068 31052 12078 31108
rect 5506 30940 5516 30996
rect 5572 30940 5582 30996
rect 11330 30940 11340 30996
rect 11396 30940 12124 30996
rect 12180 30940 12190 30996
rect 15092 30940 36988 30996
rect 37044 30940 37054 30996
rect 5516 30884 5572 30940
rect 15092 30884 15148 30940
rect 2258 30828 2268 30884
rect 2324 30828 4732 30884
rect 4788 30828 5180 30884
rect 5236 30828 5246 30884
rect 5516 30828 5964 30884
rect 6020 30828 6300 30884
rect 6356 30828 15148 30884
rect 25330 30828 25340 30884
rect 25396 30828 28700 30884
rect 28756 30828 28766 30884
rect 40114 30828 40124 30884
rect 40180 30828 41580 30884
rect 41636 30828 57596 30884
rect 57652 30828 57662 30884
rect 9426 30604 9436 30660
rect 9492 30604 9996 30660
rect 10052 30604 10062 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 5954 30492 5964 30548
rect 6020 30492 6524 30548
rect 6580 30492 8540 30548
rect 8596 30492 8606 30548
rect 9650 30492 9660 30548
rect 9716 30492 10444 30548
rect 10500 30492 10510 30548
rect 17490 30492 17500 30548
rect 17556 30492 17948 30548
rect 18004 30492 18014 30548
rect 5506 30380 5516 30436
rect 5572 30380 9212 30436
rect 9268 30380 9278 30436
rect 9426 30380 9436 30436
rect 9492 30380 11788 30436
rect 11844 30380 11854 30436
rect 18050 30380 18060 30436
rect 18116 30380 19180 30436
rect 19236 30380 19246 30436
rect 2146 30268 2156 30324
rect 2212 30268 5740 30324
rect 5796 30268 5806 30324
rect 6066 30268 6076 30324
rect 6132 30268 17052 30324
rect 17108 30268 17724 30324
rect 17780 30268 17790 30324
rect 41010 30268 41020 30324
rect 41076 30268 41412 30324
rect 41356 30212 41412 30268
rect 9874 30156 9884 30212
rect 9940 30156 12348 30212
rect 12404 30156 13132 30212
rect 13188 30156 13198 30212
rect 16034 30156 16044 30212
rect 16100 30156 17164 30212
rect 17220 30156 17836 30212
rect 17892 30156 18620 30212
rect 18676 30156 18686 30212
rect 19618 30156 19628 30212
rect 19684 30156 21644 30212
rect 21700 30156 26124 30212
rect 26180 30156 26190 30212
rect 33618 30156 33628 30212
rect 33684 30156 37436 30212
rect 37492 30156 37996 30212
rect 38052 30156 38062 30212
rect 41346 30156 41356 30212
rect 41412 30156 41422 30212
rect 10098 30044 10108 30100
rect 10164 30044 10332 30100
rect 10388 30044 10668 30100
rect 10724 30044 10734 30100
rect 12226 30044 12236 30100
rect 12292 30044 12796 30100
rect 12852 30044 12862 30100
rect 13794 30044 13804 30100
rect 13860 30044 14364 30100
rect 14420 30044 14430 30100
rect 14914 30044 14924 30100
rect 14980 30044 15484 30100
rect 15540 30044 18788 30100
rect 18946 30044 18956 30100
rect 19012 30044 19964 30100
rect 20020 30044 20030 30100
rect 20402 30044 20412 30100
rect 20468 30044 20860 30100
rect 20916 30044 22764 30100
rect 22820 30044 26908 30100
rect 26964 30044 28028 30100
rect 28084 30044 28094 30100
rect 18732 29988 18788 30044
rect 11330 29932 11340 29988
rect 11396 29932 12572 29988
rect 12628 29932 12638 29988
rect 13234 29932 13244 29988
rect 13300 29932 18508 29988
rect 18564 29932 18574 29988
rect 18732 29932 22092 29988
rect 22148 29932 22158 29988
rect 31602 29932 31612 29988
rect 31668 29932 32172 29988
rect 32228 29932 32238 29988
rect 16818 29820 16828 29876
rect 16884 29820 18284 29876
rect 18340 29820 18350 29876
rect 20402 29820 20412 29876
rect 20468 29820 21868 29876
rect 21924 29820 22316 29876
rect 22372 29820 22382 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 200 29652 800 29736
rect 22082 29708 22092 29764
rect 22148 29708 24948 29764
rect 24892 29652 24948 29708
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 10994 29596 11004 29652
rect 11060 29596 11116 29652
rect 11172 29596 11182 29652
rect 18386 29596 18396 29652
rect 18452 29596 19068 29652
rect 19124 29596 22204 29652
rect 22260 29596 22270 29652
rect 24882 29596 24892 29652
rect 24948 29596 25676 29652
rect 25732 29596 25742 29652
rect 200 29512 800 29596
rect 9650 29484 9660 29540
rect 9716 29484 12236 29540
rect 12292 29484 12302 29540
rect 18274 29484 18284 29540
rect 18340 29484 19516 29540
rect 19572 29484 20860 29540
rect 20916 29484 20926 29540
rect 23538 29484 23548 29540
rect 23604 29484 23642 29540
rect 10546 29372 10556 29428
rect 10612 29372 11340 29428
rect 11396 29372 11406 29428
rect 9314 29260 9324 29316
rect 9380 29260 11340 29316
rect 11396 29260 15484 29316
rect 15540 29260 15550 29316
rect 28914 29260 28924 29316
rect 28980 29260 32172 29316
rect 32228 29260 32732 29316
rect 32788 29260 32798 29316
rect 34514 29260 34524 29316
rect 34580 29260 35756 29316
rect 35812 29260 35822 29316
rect 11078 29148 11116 29204
rect 11172 29148 11182 29204
rect 28466 29148 28476 29204
rect 28532 29148 38108 29204
rect 38164 29148 38174 29204
rect 23090 29036 23100 29092
rect 23156 29036 23436 29092
rect 23492 29036 23502 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 25666 28924 25676 28980
rect 25732 28924 26460 28980
rect 26516 28924 34636 28980
rect 34692 28924 34702 28980
rect 35746 28924 35756 28980
rect 35812 28924 36764 28980
rect 36820 28924 36830 28980
rect 59200 28868 59800 29064
rect 12338 28812 12348 28868
rect 12404 28812 12908 28868
rect 12964 28812 13916 28868
rect 13972 28812 13982 28868
rect 17938 28812 17948 28868
rect 18004 28812 23324 28868
rect 23380 28812 23390 28868
rect 24210 28812 24220 28868
rect 24276 28812 24286 28868
rect 28018 28812 28028 28868
rect 28084 28812 33292 28868
rect 33348 28812 33628 28868
rect 33684 28812 33694 28868
rect 35298 28812 35308 28868
rect 35364 28812 39340 28868
rect 39396 28812 39406 28868
rect 58146 28812 58156 28868
rect 58212 28840 59800 28868
rect 58212 28812 59304 28840
rect 12562 28700 12572 28756
rect 12628 28700 13580 28756
rect 13636 28700 13646 28756
rect 16930 28700 16940 28756
rect 16996 28700 18508 28756
rect 18564 28700 18732 28756
rect 18788 28700 18798 28756
rect 24220 28644 24276 28812
rect 26450 28700 26460 28756
rect 26516 28700 26908 28756
rect 26964 28700 27468 28756
rect 27524 28700 27534 28756
rect 27906 28700 27916 28756
rect 27972 28700 28476 28756
rect 28532 28700 28542 28756
rect 28802 28700 28812 28756
rect 28868 28700 32620 28756
rect 32676 28700 33740 28756
rect 33796 28700 33806 28756
rect 34626 28700 34636 28756
rect 34692 28700 35532 28756
rect 35588 28700 37660 28756
rect 37716 28700 37726 28756
rect 10546 28588 10556 28644
rect 10612 28588 12012 28644
rect 12068 28588 12078 28644
rect 16594 28588 16604 28644
rect 16660 28588 17780 28644
rect 18162 28588 18172 28644
rect 18228 28588 23100 28644
rect 23156 28588 23166 28644
rect 23426 28588 23436 28644
rect 23492 28588 24668 28644
rect 24724 28588 25228 28644
rect 25284 28588 28028 28644
rect 28084 28588 28094 28644
rect 32834 28588 32844 28644
rect 32900 28588 35308 28644
rect 35364 28588 35374 28644
rect 38098 28588 38108 28644
rect 38164 28588 39564 28644
rect 39620 28588 39630 28644
rect 39890 28588 39900 28644
rect 39956 28588 40460 28644
rect 40516 28588 41244 28644
rect 41300 28588 41310 28644
rect 17724 28532 17780 28588
rect 17714 28476 17724 28532
rect 17780 28476 17790 28532
rect 23538 28476 23548 28532
rect 23604 28476 24220 28532
rect 24276 28476 28588 28532
rect 28644 28476 28654 28532
rect 29250 28476 29260 28532
rect 29316 28476 31164 28532
rect 31220 28476 32396 28532
rect 32452 28476 32462 28532
rect 12450 28364 12460 28420
rect 12516 28364 35420 28420
rect 35476 28364 35486 28420
rect 41682 28364 41692 28420
rect 41748 28364 42252 28420
rect 42308 28364 42318 28420
rect 34066 28252 34076 28308
rect 34132 28252 36316 28308
rect 36372 28252 38556 28308
rect 38612 28252 39116 28308
rect 39172 28252 39182 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 6066 28028 6076 28084
rect 6132 28028 6300 28084
rect 6356 28028 7308 28084
rect 7364 28028 7374 28084
rect 22418 28028 22428 28084
rect 22484 28028 28700 28084
rect 28756 28028 29260 28084
rect 29316 28028 29326 28084
rect 23762 27916 23772 27972
rect 23828 27916 24108 27972
rect 24164 27916 24174 27972
rect 6290 27804 6300 27860
rect 6356 27804 6748 27860
rect 6804 27804 6814 27860
rect 10322 27804 10332 27860
rect 10388 27804 11004 27860
rect 11060 27804 11564 27860
rect 11620 27804 11630 27860
rect 19506 27804 19516 27860
rect 19572 27804 25900 27860
rect 25956 27804 25966 27860
rect 6066 27692 6076 27748
rect 6132 27692 10108 27748
rect 10164 27692 10174 27748
rect 20178 27692 20188 27748
rect 20244 27692 20524 27748
rect 20580 27692 27916 27748
rect 27972 27692 27982 27748
rect 32722 27692 32732 27748
rect 32788 27692 36092 27748
rect 36148 27692 56252 27748
rect 56308 27692 56318 27748
rect 10322 27580 10332 27636
rect 10388 27580 11452 27636
rect 11508 27580 11518 27636
rect 21970 27580 21980 27636
rect 22036 27580 23548 27636
rect 23604 27580 24668 27636
rect 24724 27580 28700 27636
rect 28756 27580 28766 27636
rect 23314 27468 23324 27524
rect 23380 27468 23996 27524
rect 24052 27468 27132 27524
rect 27188 27468 27198 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 23426 27356 23436 27412
rect 23492 27356 25116 27412
rect 25172 27356 25182 27412
rect 7634 27244 7644 27300
rect 7700 27244 15148 27300
rect 15092 27076 15148 27244
rect 19180 27244 21924 27300
rect 22306 27244 22316 27300
rect 22372 27244 26012 27300
rect 26068 27244 27020 27300
rect 27076 27244 27086 27300
rect 28578 27244 28588 27300
rect 28644 27244 29484 27300
rect 29540 27244 33964 27300
rect 34020 27244 34030 27300
rect 19180 27188 19236 27244
rect 21868 27188 21924 27244
rect 18274 27132 18284 27188
rect 18340 27132 19180 27188
rect 19236 27132 19246 27188
rect 19394 27132 19404 27188
rect 19460 27132 20188 27188
rect 20244 27132 20254 27188
rect 21858 27132 21868 27188
rect 21924 27132 22428 27188
rect 22484 27132 22494 27188
rect 24434 27132 24444 27188
rect 24500 27132 25676 27188
rect 25732 27132 25742 27188
rect 25890 27132 25900 27188
rect 25956 27132 26908 27188
rect 27906 27132 27916 27188
rect 27972 27132 31276 27188
rect 31332 27132 31612 27188
rect 31668 27132 33292 27188
rect 33348 27132 33358 27188
rect 11666 27020 11676 27076
rect 11732 27020 12124 27076
rect 12180 27020 12190 27076
rect 15092 27020 17388 27076
rect 17444 27020 19628 27076
rect 19684 27020 20188 27076
rect 23202 27020 23212 27076
rect 23268 27020 25116 27076
rect 25172 27020 25182 27076
rect 3042 26908 3052 26964
rect 3108 26908 3500 26964
rect 3556 26908 10556 26964
rect 10612 26908 10622 26964
rect 17826 26908 17836 26964
rect 17892 26908 19516 26964
rect 19572 26908 19582 26964
rect 20132 26852 20188 27020
rect 26852 26964 26908 27132
rect 27682 27020 27692 27076
rect 27748 27020 28252 27076
rect 28308 27020 28318 27076
rect 28690 27020 28700 27076
rect 28756 27020 31724 27076
rect 31780 27020 32732 27076
rect 32788 27020 32798 27076
rect 28700 26964 28756 27020
rect 22530 26908 22540 26964
rect 22596 26908 24668 26964
rect 24724 26908 24734 26964
rect 25218 26908 25228 26964
rect 25284 26908 26460 26964
rect 26516 26908 26526 26964
rect 26852 26908 28756 26964
rect 35970 26908 35980 26964
rect 36036 26908 42028 26964
rect 42084 26908 42094 26964
rect 20132 26796 27132 26852
rect 27188 26796 27198 26852
rect 10210 26684 10220 26740
rect 10276 26684 12012 26740
rect 12068 26684 12460 26740
rect 12516 26684 12526 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 2370 26572 2380 26628
rect 2436 26572 7756 26628
rect 7812 26572 7822 26628
rect 10220 26572 11340 26628
rect 11396 26572 11406 26628
rect 10220 26516 10276 26572
rect 10210 26460 10220 26516
rect 10276 26460 10286 26516
rect 27234 26460 27244 26516
rect 27300 26460 27804 26516
rect 27860 26460 27870 26516
rect 41906 26460 41916 26516
rect 41972 26460 42700 26516
rect 42756 26460 42766 26516
rect 728 26376 2156 26404
rect 200 26348 2156 26376
rect 2212 26348 2222 26404
rect 39890 26348 39900 26404
rect 39956 26348 41580 26404
rect 41636 26348 41646 26404
rect 200 26152 800 26348
rect 4274 26012 4284 26068
rect 4340 26012 10220 26068
rect 10276 26012 10286 26068
rect 10882 26012 10892 26068
rect 10948 26012 11900 26068
rect 11956 26012 11966 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 59200 25620 59800 25704
rect 22418 25564 22428 25620
rect 22484 25564 22988 25620
rect 23044 25564 24108 25620
rect 24164 25564 24174 25620
rect 57810 25564 57820 25620
rect 57876 25564 59800 25620
rect 59200 25480 59800 25564
rect 9762 25340 9772 25396
rect 9828 25340 10332 25396
rect 10388 25340 10398 25396
rect 19618 25228 19628 25284
rect 19684 25228 22876 25284
rect 22932 25228 22942 25284
rect 24098 25228 24108 25284
rect 24164 25228 24174 25284
rect 24108 25172 24164 25228
rect 23650 25116 23660 25172
rect 23716 25116 24668 25172
rect 24724 25116 24734 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 24098 25004 24108 25060
rect 24164 25004 24332 25060
rect 24388 25004 24398 25060
rect 26898 25004 26908 25060
rect 26964 25004 27132 25060
rect 27188 25004 28364 25060
rect 28420 25004 28924 25060
rect 28980 25004 28990 25060
rect 23538 24892 23548 24948
rect 23604 24892 24332 24948
rect 24388 24892 24668 24948
rect 24724 24892 24734 24948
rect 27458 24892 27468 24948
rect 27524 24892 28588 24948
rect 28644 24892 28654 24948
rect 10546 24780 10556 24836
rect 10612 24780 11340 24836
rect 11396 24780 12236 24836
rect 12292 24780 12302 24836
rect 18162 24780 18172 24836
rect 18228 24780 22428 24836
rect 22484 24780 22494 24836
rect 27906 24780 27916 24836
rect 27972 24780 28812 24836
rect 28868 24780 28878 24836
rect 11106 24668 11116 24724
rect 11172 24668 11788 24724
rect 11844 24668 11854 24724
rect 23986 24668 23996 24724
rect 24052 24668 24220 24724
rect 24276 24668 24286 24724
rect 18050 24556 18060 24612
rect 18116 24556 19628 24612
rect 19684 24556 19694 24612
rect 21858 24556 21868 24612
rect 21924 24556 22428 24612
rect 22484 24556 22494 24612
rect 22754 24556 22764 24612
rect 22820 24556 23660 24612
rect 23716 24556 24444 24612
rect 24500 24556 24510 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 24322 24108 24332 24164
rect 24388 24108 26348 24164
rect 26404 24108 26414 24164
rect 26348 24052 26404 24108
rect 3042 23996 3052 24052
rect 3108 23996 3612 24052
rect 3668 23996 5852 24052
rect 5908 23996 5918 24052
rect 24210 23996 24220 24052
rect 24276 23996 24286 24052
rect 26348 23996 32508 24052
rect 32564 23996 32574 24052
rect 24220 23828 24276 23996
rect 17714 23772 17724 23828
rect 17780 23772 22316 23828
rect 22372 23772 23212 23828
rect 23268 23772 24276 23828
rect 728 23688 2156 23716
rect 200 23660 2156 23688
rect 2212 23660 2222 23716
rect 3490 23660 3500 23716
rect 3556 23660 6860 23716
rect 6916 23660 21196 23716
rect 21252 23660 21644 23716
rect 21700 23660 23100 23716
rect 23156 23660 23548 23716
rect 23604 23660 24220 23716
rect 24276 23660 24286 23716
rect 200 23464 800 23660
rect 22978 23548 22988 23604
rect 23044 23548 23548 23604
rect 23604 23548 23614 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 10434 23436 10444 23492
rect 10500 23436 11340 23492
rect 11396 23436 17164 23492
rect 17220 23436 17948 23492
rect 18004 23436 18620 23492
rect 18676 23436 19180 23492
rect 19236 23436 19246 23492
rect 17378 23324 17388 23380
rect 17444 23324 17836 23380
rect 17892 23324 18172 23380
rect 18228 23324 18844 23380
rect 18900 23324 18910 23380
rect 46722 23212 46732 23268
rect 46788 23212 57708 23268
rect 57764 23212 57774 23268
rect 10658 22988 10668 23044
rect 10724 22988 11004 23044
rect 11060 22988 11676 23044
rect 11732 22988 16940 23044
rect 16996 22988 18396 23044
rect 18452 22988 21644 23044
rect 21700 22988 21980 23044
rect 22036 22988 22764 23044
rect 22820 22988 22830 23044
rect 58034 22988 58044 23044
rect 58100 23016 59304 23044
rect 58100 22988 59800 23016
rect 59200 22792 59800 22988
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 3602 22316 3612 22372
rect 3668 22316 10332 22372
rect 10388 22316 11676 22372
rect 11732 22316 12236 22372
rect 12292 22316 12302 22372
rect 9986 22204 9996 22260
rect 10052 22204 11788 22260
rect 11844 22204 11854 22260
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 3938 21756 3948 21812
rect 4004 21756 9436 21812
rect 9492 21756 9502 21812
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 728 21000 2044 21028
rect 200 20972 2044 21000
rect 2100 20972 2110 21028
rect 200 20776 800 20972
rect 46498 20636 46508 20692
rect 46564 20636 57708 20692
rect 57764 20636 57774 20692
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 57250 20300 57260 20356
rect 57316 20300 58044 20356
rect 58100 20328 59304 20356
rect 58100 20300 59800 20328
rect 59200 20104 59800 20300
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 2146 18620 2156 18676
rect 2212 18620 3724 18676
rect 3780 18620 3790 18676
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 200 17556 800 17640
rect 200 17500 1820 17556
rect 1876 17500 1886 17556
rect 41122 17500 41132 17556
rect 41188 17500 57708 17556
rect 57764 17500 57774 17556
rect 200 17416 800 17500
rect 57250 17388 57260 17444
rect 57316 17388 58044 17444
rect 58100 17388 58110 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 58034 16940 58044 16996
rect 58100 16968 59304 16996
rect 58100 16940 59800 16968
rect 59200 16744 59800 16940
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 200 14756 800 14952
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 200 14728 1820 14756
rect 728 14700 1820 14728
rect 1876 14700 1886 14756
rect 51314 14588 51324 14644
rect 51380 14588 56364 14644
rect 56420 14588 56812 14644
rect 56868 14588 56878 14644
rect 57698 14252 57708 14308
rect 57764 14280 59304 14308
rect 57764 14252 59800 14280
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 59200 14056 59800 14252
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 3042 12348 3052 12404
rect 3108 12348 3500 12404
rect 3556 12348 7532 12404
rect 7588 12348 7598 12404
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 728 11592 2044 11620
rect 200 11564 2044 11592
rect 2100 11564 2110 11620
rect 200 11368 800 11564
rect 28802 11116 28812 11172
rect 28868 11116 56364 11172
rect 56420 11116 56812 11172
rect 56868 11116 56878 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 57698 10892 57708 10948
rect 57764 10920 59304 10948
rect 57764 10892 59800 10920
rect 59200 10696 59800 10892
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 200 8708 800 8904
rect 200 8680 1820 8708
rect 728 8652 1820 8680
rect 1876 8652 1886 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 59200 8148 59800 8232
rect 40338 8092 40348 8148
rect 40404 8092 57708 8148
rect 57764 8092 57774 8148
rect 58034 8092 58044 8148
rect 58100 8092 59800 8148
rect 58044 8036 58100 8092
rect 57250 7980 57260 8036
rect 57316 7980 58100 8036
rect 59200 8008 59800 8092
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 3042 6076 3052 6132
rect 3108 6076 3500 6132
rect 3556 6076 6412 6132
rect 6468 6076 6478 6132
rect 728 5544 2044 5572
rect 200 5516 2044 5544
rect 2100 5516 2110 5572
rect 200 5320 800 5516
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 11330 5292 11340 5348
rect 11396 5292 16492 5348
rect 16548 5292 16558 5348
rect 3042 5180 3052 5236
rect 3108 5180 3612 5236
rect 3668 5180 6188 5236
rect 6244 5180 6254 5236
rect 58034 5180 58044 5236
rect 58100 5180 59332 5236
rect 59276 5012 59332 5180
rect 802 4956 812 5012
rect 868 4956 2156 5012
rect 2212 4956 2222 5012
rect 57250 4956 57260 5012
rect 57316 4956 58044 5012
rect 58100 4956 58110 5012
rect 59164 4956 59332 5012
rect 59164 4900 59220 4956
rect 59164 4872 59304 4900
rect 59164 4844 59800 4872
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 59200 4648 59800 4844
rect 11106 4508 11116 4564
rect 11172 4508 12348 4564
rect 12404 4508 12414 4564
rect 56802 4172 56812 4228
rect 56868 4172 58044 4228
rect 58100 4172 58110 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 11778 3612 11788 3668
rect 11844 3612 16828 3668
rect 16884 3612 17724 3668
rect 17780 3612 17790 3668
rect 44258 3612 44268 3668
rect 44324 3612 45612 3668
rect 45668 3612 45678 3668
rect 42466 3500 42476 3556
rect 42532 3500 56028 3556
rect 56084 3500 56700 3556
rect 56756 3500 56766 3556
rect 8866 3388 8876 3444
rect 8932 3388 9996 3444
rect 10052 3388 10062 3444
rect 20738 3388 20748 3444
rect 20804 3388 21420 3444
rect 21476 3388 21486 3444
rect 32386 3388 32396 3444
rect 32452 3388 34076 3444
rect 34132 3388 34142 3444
rect 48178 3388 48188 3444
rect 48244 3388 49196 3444
rect 49252 3388 49262 3444
rect 50418 3388 50428 3444
rect 50484 3388 50988 3444
rect 51044 3388 51054 3444
rect 56578 3388 56588 3444
rect 56644 3388 57596 3444
rect 57652 3388 57662 3444
rect 21746 3276 21756 3332
rect 21812 3276 28140 3332
rect 28196 3276 28206 3332
rect 30146 3276 30156 3332
rect 30212 3276 31612 3332
rect 31668 3276 31678 3332
rect 42354 3276 42364 3332
rect 42420 3276 50652 3332
rect 50708 3276 50718 3332
rect 40674 3164 40684 3220
rect 40740 3164 48860 3220
rect 48916 3164 48926 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 728 2856 2044 2884
rect 200 2828 2044 2856
rect 2100 2828 2110 2884
rect 58034 2828 58044 2884
rect 58100 2828 59332 2884
rect 200 2632 800 2828
rect 59276 2324 59332 2828
rect 59164 2268 59332 2324
rect 59164 2212 59220 2268
rect 59164 2184 59304 2212
rect 59164 2156 59800 2184
rect 59200 1960 59800 2156
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 24108 46284 24164 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 24108 46060 24164 46116
rect 32620 45724 32676 45780
rect 30716 45500 30772 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 31164 45500 31220 45556
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 17388 45276 17444 45332
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4844 39004 4900 39060
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 4844 38332 4900 38388
rect 39452 37772 39508 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 19068 37436 19124 37492
rect 32620 37436 32676 37492
rect 19180 37212 19236 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 35644 36764 35700 36820
rect 32732 36652 32788 36708
rect 17388 36540 17444 36596
rect 19068 36540 19124 36596
rect 32844 36204 32900 36260
rect 19180 36092 19236 36148
rect 35644 36092 35700 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 29148 35196 29204 35252
rect 39452 34972 39508 35028
rect 29148 34860 29204 34916
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 26796 33628 26852 33684
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 26796 32956 26852 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 24332 31500 24388 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 11116 29596 11172 29652
rect 23548 29484 23604 29540
rect 11340 29260 11396 29316
rect 11116 29148 11172 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 25900 27804 25956 27860
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 25900 27132 25956 27188
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 11340 26572 11396 26628
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 24108 25564 24164 25620
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 24332 25004 24388 25060
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 23548 23660 23604 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 17388 45332 17444 45342
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4844 39060 4900 39070
rect 4844 38388 4900 39004
rect 4844 38322 4900 38332
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 17388 36596 17444 45276
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 17388 36530 17444 36540
rect 19068 37492 19124 37502
rect 19068 36596 19124 37436
rect 19068 36530 19124 36540
rect 19180 37268 19236 37278
rect 19180 36148 19236 37212
rect 19180 36082 19236 36092
rect 19808 36092 20128 37604
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 11116 29652 11172 29662
rect 11116 29204 11172 29596
rect 11116 29138 11172 29148
rect 11340 29316 11396 29326
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 11340 26628 11396 29260
rect 11340 26562 11396 26572
rect 19808 28252 20128 29764
rect 24108 46340 24164 46350
rect 24108 46116 24164 46284
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 23548 29540 23604 29550
rect 23548 23716 23604 29484
rect 24108 25620 24164 46060
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 32620 45780 32676 45790
rect 30716 45556 30772 45566
rect 31164 45556 31220 45566
rect 30772 45500 31164 45556
rect 30716 45490 30772 45500
rect 31164 45490 31220 45500
rect 32620 37492 32676 45724
rect 32620 37426 32676 37436
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 39452 37828 39508 37838
rect 32732 36708 32788 36718
rect 32788 36652 32900 36708
rect 32732 36642 32788 36652
rect 32844 36260 32900 36652
rect 32844 36194 32900 36204
rect 35168 35308 35488 36820
rect 35644 36820 35700 36830
rect 35644 36148 35700 36764
rect 35644 36082 35700 36092
rect 29148 35252 29204 35262
rect 29148 34916 29204 35196
rect 29148 34850 29204 34860
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 39452 35028 39508 37772
rect 39452 34962 39508 34972
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 26796 33684 26852 33694
rect 26796 33012 26852 33628
rect 26796 32946 26852 32956
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 24108 25554 24164 25564
rect 24332 31556 24388 31566
rect 24332 25060 24388 31500
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 25900 27860 25956 27870
rect 25900 27188 25956 27804
rect 25900 27122 25956 27132
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 24332 24994 24388 25004
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 23548 23650 23604 23660
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A1 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 17696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A2
timestamp 1666464484
transform 1 0 19376 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A1
timestamp 1666464484
transform 1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A2
timestamp 1666464484
transform 1 0 18144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A1
timestamp 1666464484
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A2
timestamp 1666464484
transform 1 0 26320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A3
timestamp 1666464484
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__I
timestamp 1666464484
transform 1 0 42448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I
timestamp 1666464484
transform 1 0 38864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A1
timestamp 1666464484
transform -1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A2
timestamp 1666464484
transform 1 0 34048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__A1
timestamp 1666464484
transform -1 0 37632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__A2
timestamp 1666464484
transform 1 0 37856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__A3
timestamp 1666464484
transform -1 0 36512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__A4
timestamp 1666464484
transform 1 0 37408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A1
timestamp 1666464484
transform 1 0 35616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A3
timestamp 1666464484
transform 1 0 36064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A4
timestamp 1666464484
transform 1 0 36512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A2
timestamp 1666464484
transform 1 0 24640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A3
timestamp 1666464484
transform 1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A1
timestamp 1666464484
transform 1 0 24080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A2
timestamp 1666464484
transform 1 0 24528 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A3
timestamp 1666464484
transform 1 0 27328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A4
timestamp 1666464484
transform 1 0 24976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__I
timestamp 1666464484
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A1
timestamp 1666464484
transform 1 0 47264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A2
timestamp 1666464484
transform 1 0 49056 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__B
timestamp 1666464484
transform 1 0 46816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A1
timestamp 1666464484
transform 1 0 46592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A2
timestamp 1666464484
transform 1 0 47040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A3
timestamp 1666464484
transform 1 0 47488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__A1
timestamp 1666464484
transform -1 0 48832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__A1
timestamp 1666464484
transform -1 0 40768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A1
timestamp 1666464484
transform 1 0 39424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A2
timestamp 1666464484
transform -1 0 41664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__B1
timestamp 1666464484
transform 1 0 38976 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__B2
timestamp 1666464484
transform 1 0 38528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A1
timestamp 1666464484
transform 1 0 52640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A2
timestamp 1666464484
transform 1 0 53088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__A1
timestamp 1666464484
transform 1 0 52192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__A1
timestamp 1666464484
transform 1 0 39424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__A2
timestamp 1666464484
transform -1 0 38528 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__I
timestamp 1666464484
transform 1 0 46032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__A1
timestamp 1666464484
transform 1 0 41440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__A2
timestamp 1666464484
transform 1 0 42784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__B2
timestamp 1666464484
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__I
timestamp 1666464484
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A1
timestamp 1666464484
transform 1 0 13664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A2
timestamp 1666464484
transform 1 0 14672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A3
timestamp 1666464484
transform 1 0 15568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__277__A1
timestamp 1666464484
transform 1 0 12320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A1
timestamp 1666464484
transform 1 0 5936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A2
timestamp 1666464484
transform -1 0 4816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__A1
timestamp 1666464484
transform 1 0 10416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__B2
timestamp 1666464484
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__I
timestamp 1666464484
transform 1 0 11312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I
timestamp 1666464484
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A1
timestamp 1666464484
transform 1 0 30464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A2
timestamp 1666464484
transform 1 0 30016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1666464484
transform 1 0 35504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A1
timestamp 1666464484
transform 1 0 40656 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A2
timestamp 1666464484
transform 1 0 41440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__A1
timestamp 1666464484
transform 1 0 35952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__B2
timestamp 1666464484
transform 1 0 36176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A1
timestamp 1666464484
transform 1 0 26320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A2
timestamp 1666464484
transform 1 0 25872 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A3
timestamp 1666464484
transform 1 0 26320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A4
timestamp 1666464484
transform 1 0 26768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__A1
timestamp 1666464484
transform 1 0 42448 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__A2
timestamp 1666464484
transform -1 0 42224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A1
timestamp 1666464484
transform 1 0 40880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A1
timestamp 1666464484
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1666464484
transform -1 0 41664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__A1
timestamp 1666464484
transform -1 0 37184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__B1
timestamp 1666464484
transform 1 0 38976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__B2
timestamp 1666464484
transform 1 0 37408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A1
timestamp 1666464484
transform 1 0 17584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A2
timestamp 1666464484
transform 1 0 19488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A1
timestamp 1666464484
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A2
timestamp 1666464484
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A3
timestamp 1666464484
transform 1 0 21616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__I
timestamp 1666464484
transform 1 0 51296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1666464484
transform 1 0 46032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A1
timestamp 1666464484
transform 1 0 35728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A2
timestamp 1666464484
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A3
timestamp 1666464484
transform -1 0 35056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A4
timestamp 1666464484
transform -1 0 35504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A1
timestamp 1666464484
transform 1 0 41888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A2
timestamp 1666464484
transform 1 0 41552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A3
timestamp 1666464484
transform -1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A1
timestamp 1666464484
transform 1 0 23968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A2
timestamp 1666464484
transform -1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A3
timestamp 1666464484
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A4
timestamp 1666464484
transform 1 0 26544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A1
timestamp 1666464484
transform 1 0 27216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A2
timestamp 1666464484
transform -1 0 27888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__B
timestamp 1666464484
transform 1 0 26768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A1
timestamp 1666464484
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A1
timestamp 1666464484
transform 1 0 32592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A1
timestamp 1666464484
transform -1 0 9072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A2
timestamp 1666464484
transform 1 0 7728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A1
timestamp 1666464484
transform 1 0 18480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A2
timestamp 1666464484
transform 1 0 20496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A3
timestamp 1666464484
transform -1 0 19152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__B1
timestamp 1666464484
transform 1 0 20944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__B2
timestamp 1666464484
transform 1 0 18480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A1
timestamp 1666464484
transform 1 0 33936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1666464484
transform 1 0 34384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__A1
timestamp 1666464484
transform 1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__A2
timestamp 1666464484
transform 1 0 24304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1666464484
transform 1 0 14896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__A1
timestamp 1666464484
transform 1 0 24192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__A2
timestamp 1666464484
transform -1 0 26432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__B1
timestamp 1666464484
transform 1 0 26656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__B2
timestamp 1666464484
transform 1 0 23744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A1
timestamp 1666464484
transform 1 0 13328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A2
timestamp 1666464484
transform 1 0 14896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A1
timestamp 1666464484
transform 1 0 13104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A1
timestamp 1666464484
transform 1 0 5152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__A1
timestamp 1666464484
transform -1 0 11536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__A3
timestamp 1666464484
transform 1 0 10864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__B1
timestamp 1666464484
transform 1 0 15344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__B2
timestamp 1666464484
transform 1 0 14448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1666464484
transform 1 0 16912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A1
timestamp 1666464484
transform 1 0 20832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A3
timestamp 1666464484
transform 1 0 20384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A4
timestamp 1666464484
transform -1 0 21728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A1
timestamp 1666464484
transform 1 0 16016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A2
timestamp 1666464484
transform 1 0 17472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A3
timestamp 1666464484
transform -1 0 18144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__A1
timestamp 1666464484
transform 1 0 19824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__A1
timestamp 1666464484
transform 1 0 37744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__A2
timestamp 1666464484
transform 1 0 38192 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A1
timestamp 1666464484
transform 1 0 18256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A3
timestamp 1666464484
transform -1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__B2
timestamp 1666464484
transform 1 0 17808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1666464484
transform 1 0 16464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A1
timestamp 1666464484
transform 1 0 14336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A2
timestamp 1666464484
transform 1 0 14112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__A1
timestamp 1666464484
transform 1 0 15344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__A1
timestamp 1666464484
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__A2
timestamp 1666464484
transform -1 0 35504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__A1
timestamp 1666464484
transform 1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__A3
timestamp 1666464484
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__B2
timestamp 1666464484
transform 1 0 16912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A1
timestamp 1666464484
transform 1 0 13552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A2
timestamp 1666464484
transform -1 0 12992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__B
timestamp 1666464484
transform 1 0 13104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__A1
timestamp 1666464484
transform 1 0 4480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1666464484
transform 1 0 14672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A1
timestamp 1666464484
transform 1 0 12880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A3
timestamp 1666464484
transform -1 0 11536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__B2
timestamp 1666464484
transform 1 0 14000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__I
timestamp 1666464484
transform 1 0 21728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A1
timestamp 1666464484
transform 1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A2
timestamp 1666464484
transform -1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A3
timestamp 1666464484
transform 1 0 27776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A1
timestamp 1666464484
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A3
timestamp 1666464484
transform 1 0 26432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A4
timestamp 1666464484
transform 1 0 29456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A1
timestamp 1666464484
transform 1 0 26432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A2
timestamp 1666464484
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__A1
timestamp 1666464484
transform 1 0 27776 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__A1
timestamp 1666464484
transform 1 0 31696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__A2
timestamp 1666464484
transform 1 0 31248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__I
timestamp 1666464484
transform 1 0 28224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__A1
timestamp 1666464484
transform -1 0 26992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__B2
timestamp 1666464484
transform 1 0 28560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__I
timestamp 1666464484
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__I
timestamp 1666464484
transform 1 0 32144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A1
timestamp 1666464484
transform 1 0 33264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A2
timestamp 1666464484
transform 1 0 34384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A1
timestamp 1666464484
transform 1 0 31696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A2
timestamp 1666464484
transform 1 0 31248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A3
timestamp 1666464484
transform 1 0 32144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A2
timestamp 1666464484
transform 1 0 38528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__B
timestamp 1666464484
transform 1 0 38080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__C
timestamp 1666464484
transform -1 0 40544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__A1
timestamp 1666464484
transform -1 0 42784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__A2
timestamp 1666464484
transform 1 0 43008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A1
timestamp 1666464484
transform 1 0 34608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__B1
timestamp 1666464484
transform 1 0 34160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__I
timestamp 1666464484
transform 1 0 36176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__A1
timestamp 1666464484
transform 1 0 31584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__A2
timestamp 1666464484
transform 1 0 31136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__A1
timestamp 1666464484
transform -1 0 35840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__A2
timestamp 1666464484
transform 1 0 35840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__A1
timestamp 1666464484
transform 1 0 36288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__B
timestamp 1666464484
transform 1 0 36960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A1
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A2
timestamp 1666464484
transform -1 0 41664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A1
timestamp 1666464484
transform 1 0 39088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__B1
timestamp 1666464484
transform 1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__B2
timestamp 1666464484
transform 1 0 38192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1666464484
transform 1 0 16128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1666464484
transform 1 0 20384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A1
timestamp 1666464484
transform 1 0 29232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__A2
timestamp 1666464484
transform 1 0 21952 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1666464484
transform 1 0 50288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A1
timestamp 1666464484
transform 1 0 23744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__B
timestamp 1666464484
transform 1 0 23296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__A1
timestamp 1666464484
transform 1 0 4480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__A1
timestamp 1666464484
transform 1 0 18256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__A3
timestamp 1666464484
transform 1 0 17808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__B2
timestamp 1666464484
transform 1 0 18704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1666464484
transform 1 0 24192 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A2
timestamp 1666464484
transform 1 0 23744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__B
timestamp 1666464484
transform 1 0 22176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__B
timestamp 1666464484
transform 1 0 24192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A1
timestamp 1666464484
transform 1 0 6496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A1
timestamp 1666464484
transform -1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A3
timestamp 1666464484
transform -1 0 17136 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__B1
timestamp 1666464484
transform -1 0 19152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__B2
timestamp 1666464484
transform 1 0 17136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A1
timestamp 1666464484
transform 1 0 33488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A2
timestamp 1666464484
transform 1 0 34832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1666464484
transform 1 0 32816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A2
timestamp 1666464484
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A3
timestamp 1666464484
transform 1 0 33264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A1
timestamp 1666464484
transform -1 0 41664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A2
timestamp 1666464484
transform 1 0 41664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A1
timestamp 1666464484
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A1
timestamp 1666464484
transform 1 0 42896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A2
timestamp 1666464484
transform -1 0 43568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__A1
timestamp 1666464484
transform 1 0 39984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__B1
timestamp 1666464484
transform 1 0 41776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__B2
timestamp 1666464484
transform 1 0 39536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__I
timestamp 1666464484
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1666464484
transform 1 0 32368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A2
timestamp 1666464484
transform 1 0 32592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__A1
timestamp 1666464484
transform 1 0 31920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__B
timestamp 1666464484
transform 1 0 30912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A1
timestamp 1666464484
transform 1 0 38976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A2
timestamp 1666464484
transform -1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A1
timestamp 1666464484
transform 1 0 29680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A3
timestamp 1666464484
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__B2
timestamp 1666464484
transform 1 0 29680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__I
timestamp 1666464484
transform -1 0 33040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A1
timestamp 1666464484
transform 1 0 36288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__A1
timestamp 1666464484
transform 1 0 34160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__B
timestamp 1666464484
transform 1 0 32256 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A1
timestamp 1666464484
transform -1 0 28336 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__A1
timestamp 1666464484
transform 1 0 28672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__A3
timestamp 1666464484
transform -1 0 27664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__B1
timestamp 1666464484
transform 1 0 30688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__B2
timestamp 1666464484
transform 1 0 27888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1666464484
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A2
timestamp 1666464484
transform 1 0 35616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__B
timestamp 1666464484
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A1
timestamp 1666464484
transform 1 0 39872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2
timestamp 1666464484
transform 1 0 40320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__A1
timestamp 1666464484
transform 1 0 37408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__B2
timestamp 1666464484
transform 1 0 37856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1666464484
transform 1 0 42000 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A2
timestamp 1666464484
transform 1 0 43120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A3
timestamp 1666464484
transform 1 0 42448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__A1
timestamp 1666464484
transform 1 0 46704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A1
timestamp 1666464484
transform 1 0 50960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1666464484
transform 1 0 49952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A1
timestamp 1666464484
transform 1 0 45136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1666464484
transform -1 0 46704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__A1
timestamp 1666464484
transform 1 0 45136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__B1
timestamp 1666464484
transform -1 0 47376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__B2
timestamp 1666464484
transform 1 0 44688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A1
timestamp 1666464484
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__B
timestamp 1666464484
transform 1 0 49392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1666464484
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A2
timestamp 1666464484
transform 1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A1
timestamp 1666464484
transform 1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__B1
timestamp 1666464484
transform 1 0 46592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__B2
timestamp 1666464484
transform 1 0 44128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__I
timestamp 1666464484
transform 1 0 40320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A1
timestamp 1666464484
transform 1 0 39872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A2
timestamp 1666464484
transform 1 0 41104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__B
timestamp 1666464484
transform -1 0 43904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A1
timestamp 1666464484
transform 1 0 43568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A2
timestamp 1666464484
transform 1 0 44912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A1
timestamp 1666464484
transform -1 0 42448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__B2
timestamp 1666464484
transform 1 0 41776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__I
timestamp 1666464484
transform 1 0 33152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__A2
timestamp 1666464484
transform 1 0 34384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__B
timestamp 1666464484
transform 1 0 39200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1666464484
transform 1 0 33040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1666464484
transform 1 0 31696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1666464484
transform 1 0 35056 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A3
timestamp 1666464484
transform -1 0 34384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__B2
timestamp 1666464484
transform 1 0 35504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I
timestamp 1666464484
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A1
timestamp 1666464484
transform 1 0 23184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A2
timestamp 1666464484
transform 1 0 23632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A1
timestamp 1666464484
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A2
timestamp 1666464484
transform -1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A2
timestamp 1666464484
transform 1 0 37408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A3
timestamp 1666464484
transform -1 0 36960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A1
timestamp 1666464484
transform 1 0 39760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A2
timestamp 1666464484
transform 1 0 42112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A1
timestamp 1666464484
transform 1 0 20832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A2
timestamp 1666464484
transform 1 0 23296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__B1
timestamp 1666464484
transform 1 0 20384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__B2
timestamp 1666464484
transform -1 0 23072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__I
timestamp 1666464484
transform 1 0 30128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A1
timestamp 1666464484
transform 1 0 24640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__A2
timestamp 1666464484
transform 1 0 26992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A1
timestamp 1666464484
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__B
timestamp 1666464484
transform 1 0 27216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1666464484
transform 1 0 42672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A2
timestamp 1666464484
transform 1 0 44016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1666464484
transform 1 0 24080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A3
timestamp 1666464484
transform -1 0 26320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__B2
timestamp 1666464484
transform 1 0 26544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1666464484
transform 1 0 19152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A2
timestamp 1666464484
transform 1 0 16912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__B
timestamp 1666464484
transform -1 0 18928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1666464484
transform 1 0 23968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__B
timestamp 1666464484
transform -1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A1
timestamp 1666464484
transform -1 0 29568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A2
timestamp 1666464484
transform -1 0 28224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1666464484
transform 1 0 22960 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A1
timestamp 1666464484
transform -1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__B2
timestamp 1666464484
transform -1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__I
timestamp 1666464484
transform -1 0 42336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1666464484
transform -1 0 36736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__I
timestamp 1666464484
transform 1 0 28672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I
timestamp 1666464484
transform 1 0 29456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__I
timestamp 1666464484
transform 1 0 31696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__I
timestamp 1666464484
transform -1 0 27888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__I
timestamp 1666464484
transform 1 0 30688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__I
timestamp 1666464484
transform 1 0 28224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__I
timestamp 1666464484
transform 1 0 27888 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1666464484
transform 1 0 29904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__I
timestamp 1666464484
transform 1 0 29120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I
timestamp 1666464484
transform -1 0 29232 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I
timestamp 1666464484
transform 1 0 37408 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1666464484
transform -1 0 26880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1666464484
transform 1 0 30016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__I
timestamp 1666464484
transform -1 0 30688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1666464484
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__I
timestamp 1666464484
transform 1 0 31136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__I
timestamp 1666464484
transform 1 0 27552 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__I
timestamp 1666464484
transform 1 0 33040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__I
timestamp 1666464484
transform 1 0 32368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__I
timestamp 1666464484
transform 1 0 32592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__I
timestamp 1666464484
transform 1 0 32368 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__I
timestamp 1666464484
transform 1 0 36848 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__I
timestamp 1666464484
transform 1 0 29456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1666464484
transform -1 0 30800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__I
timestamp 1666464484
transform 1 0 29456 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__I
timestamp 1666464484
transform 1 0 31472 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__I
timestamp 1666464484
transform 1 0 32592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__I
timestamp 1666464484
transform 1 0 31584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__I
timestamp 1666464484
transform 1 0 31920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__I
timestamp 1666464484
transform 1 0 33040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__I
timestamp 1666464484
transform 1 0 32368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__I
timestamp 1666464484
transform 1 0 32032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1666464484
transform 1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__I
timestamp 1666464484
transform 1 0 34496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__I
timestamp 1666464484
transform 1 0 50512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A1
timestamp 1666464484
transform 1 0 11760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A2
timestamp 1666464484
transform 1 0 9408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A3
timestamp 1666464484
transform 1 0 12208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A4
timestamp 1666464484
transform 1 0 11312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A1
timestamp 1666464484
transform -1 0 11424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A2
timestamp 1666464484
transform 1 0 11648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1666464484
transform -1 0 10416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A1
timestamp 1666464484
transform -1 0 9856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A2
timestamp 1666464484
transform 1 0 8176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__I
timestamp 1666464484
transform 1 0 11312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I
timestamp 1666464484
transform 1 0 41776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1666464484
transform -1 0 4704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1666464484
transform 1 0 4368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A1
timestamp 1666464484
transform 1 0 10528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A2
timestamp 1666464484
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A3
timestamp 1666464484
transform -1 0 6496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__B1
timestamp 1666464484
transform -1 0 6944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__I
timestamp 1666464484
transform 1 0 51856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__I
timestamp 1666464484
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__A1
timestamp 1666464484
transform 1 0 9744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__A2
timestamp 1666464484
transform 1 0 11760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__A3
timestamp 1666464484
transform 1 0 12208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A1
timestamp 1666464484
transform 1 0 12096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A1
timestamp 1666464484
transform -1 0 7392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1666464484
transform 1 0 6720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__I
timestamp 1666464484
transform 1 0 10192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__A1
timestamp 1666464484
transform 1 0 11984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__B2
timestamp 1666464484
transform 1 0 11536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__I
timestamp 1666464484
transform 1 0 8960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A1
timestamp 1666464484
transform 1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A2
timestamp 1666464484
transform 1 0 11312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__B
timestamp 1666464484
transform 1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A1
timestamp 1666464484
transform 1 0 35952 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A2
timestamp 1666464484
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A1
timestamp 1666464484
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A3
timestamp 1666464484
transform 1 0 11424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__B2
timestamp 1666464484
transform 1 0 11872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__I
timestamp 1666464484
transform 1 0 8512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__I
timestamp 1666464484
transform 1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__B
timestamp 1666464484
transform 1 0 11760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A1
timestamp 1666464484
transform 1 0 5488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A1
timestamp 1666464484
transform 1 0 11648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__B2
timestamp 1666464484
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A2
timestamp 1666464484
transform 1 0 10080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A1
timestamp 1666464484
transform 1 0 3136 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A2
timestamp 1666464484
transform 1 0 4480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A1
timestamp 1666464484
transform 1 0 5040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A3
timestamp 1666464484
transform 1 0 5600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__B2
timestamp 1666464484
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__I
timestamp 1666464484
transform -1 0 38640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__I
timestamp 1666464484
transform -1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__I
timestamp 1666464484
transform -1 0 27664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__I
timestamp 1666464484
transform 1 0 15120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A1
timestamp 1666464484
transform -1 0 31584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A2
timestamp 1666464484
transform 1 0 26544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A3
timestamp 1666464484
transform 1 0 26880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A4
timestamp 1666464484
transform -1 0 27216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A1
timestamp 1666464484
transform 1 0 15792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A2
timestamp 1666464484
transform -1 0 17808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A1
timestamp 1666464484
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A2
timestamp 1666464484
transform 1 0 17808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A3
timestamp 1666464484
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A4
timestamp 1666464484
transform 1 0 18256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__CLK
timestamp 1666464484
transform -1 0 19712 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__D
timestamp 1666464484
transform -1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__CLK
timestamp 1666464484
transform 1 0 19712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__D
timestamp 1666464484
transform -1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__CLK
timestamp 1666464484
transform 1 0 11200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__D
timestamp 1666464484
transform 1 0 11648 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__RN
timestamp 1666464484
transform 1 0 10752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__CLK
timestamp 1666464484
transform 1 0 19600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__D
timestamp 1666464484
transform -1 0 24304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__CLK
timestamp 1666464484
transform 1 0 11424 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__D
timestamp 1666464484
transform 1 0 11872 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__RN
timestamp 1666464484
transform -1 0 11200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__CLK
timestamp 1666464484
transform 1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__D
timestamp 1666464484
transform -1 0 23296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__RN
timestamp 1666464484
transform -1 0 23744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__CLK
timestamp 1666464484
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__D
timestamp 1666464484
transform 1 0 20384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__RN
timestamp 1666464484
transform 1 0 21504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__CLK
timestamp 1666464484
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__D
timestamp 1666464484
transform 1 0 20832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__RN
timestamp 1666464484
transform -1 0 20160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__CLK
timestamp 1666464484
transform 1 0 19824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__D
timestamp 1666464484
transform 1 0 24304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__RN
timestamp 1666464484
transform -1 0 24976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__CLK
timestamp 1666464484
transform 1 0 11872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__D
timestamp 1666464484
transform 1 0 12320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__RN
timestamp 1666464484
transform 1 0 11424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__CLK
timestamp 1666464484
transform 1 0 19600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__D
timestamp 1666464484
transform -1 0 24304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__RN
timestamp 1666464484
transform -1 0 24752 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__CLK
timestamp 1666464484
transform 1 0 12656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__D
timestamp 1666464484
transform 1 0 12432 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__RN
timestamp 1666464484
transform -1 0 12432 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__CLK
timestamp 1666464484
transform 1 0 20496 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__D
timestamp 1666464484
transform 1 0 21504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__RN
timestamp 1666464484
transform -1 0 22176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__CLK
timestamp 1666464484
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__D
timestamp 1666464484
transform 1 0 17584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__RN
timestamp 1666464484
transform 1 0 18032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__CLK
timestamp 1666464484
transform 1 0 11648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__D
timestamp 1666464484
transform 1 0 12096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__RN
timestamp 1666464484
transform -1 0 11424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__CLK
timestamp 1666464484
transform 1 0 18480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__D
timestamp 1666464484
transform -1 0 23184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__CLK
timestamp 1666464484
transform 1 0 18256 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__D
timestamp 1666464484
transform 1 0 13776 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__RN
timestamp 1666464484
transform 1 0 18704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__CLK
timestamp 1666464484
transform 1 0 9632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__D
timestamp 1666464484
transform -1 0 10864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__RN
timestamp 1666464484
transform -1 0 9856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__CLK
timestamp 1666464484
transform -1 0 11088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__D
timestamp 1666464484
transform 1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__RN
timestamp 1666464484
transform -1 0 10640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__CLK
timestamp 1666464484
transform -1 0 11088 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__D
timestamp 1666464484
transform 1 0 11312 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__RN
timestamp 1666464484
transform -1 0 10640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__CLK
timestamp 1666464484
transform 1 0 19936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__D
timestamp 1666464484
transform -1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__CLK
timestamp 1666464484
transform 1 0 19824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__D
timestamp 1666464484
transform 1 0 20272 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__RN
timestamp 1666464484
transform -1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__CLK
timestamp 1666464484
transform 1 0 18256 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__D
timestamp 1666464484
transform -1 0 23744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__CLK
timestamp 1666464484
transform 1 0 17584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__D
timestamp 1666464484
transform -1 0 18256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__RN
timestamp 1666464484
transform -1 0 18704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__CLK
timestamp 1666464484
transform 1 0 12544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__D
timestamp 1666464484
transform 1 0 12320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__RN
timestamp 1666464484
transform 1 0 12096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__CLK
timestamp 1666464484
transform 1 0 19152 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__D
timestamp 1666464484
transform -1 0 19824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__RN
timestamp 1666464484
transform 1 0 18704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__CLK
timestamp 1666464484
transform 1 0 9632 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__D
timestamp 1666464484
transform -1 0 10304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__RN
timestamp 1666464484
transform 1 0 10528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__CLK
timestamp 1666464484
transform 1 0 12096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__D
timestamp 1666464484
transform -1 0 12768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__RN
timestamp 1666464484
transform -1 0 17808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__CLK
timestamp 1666464484
transform 1 0 12208 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__D
timestamp 1666464484
transform 1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__RN
timestamp 1666464484
transform -1 0 11984 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__CLK
timestamp 1666464484
transform 1 0 10080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__D
timestamp 1666464484
transform 1 0 11200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__RN
timestamp 1666464484
transform -1 0 9856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__CLK
timestamp 1666464484
transform 1 0 10640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__D
timestamp 1666464484
transform 1 0 11088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__RN
timestamp 1666464484
transform 1 0 10192 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__CLK
timestamp 1666464484
transform 1 0 18816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__D
timestamp 1666464484
transform 1 0 14336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__RN
timestamp 1666464484
transform 1 0 19264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1666464484
transform 1 0 19376 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 15456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 21504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 15680 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 21504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 1904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform -1 0 57344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform -1 0 58240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1666464484
transform -1 0 57344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1666464484
transform -1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1666464484
transform -1 0 48272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1666464484
transform -1 0 57344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1666464484
transform -1 0 1904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1666464484
transform -1 0 1904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1666464484
transform -1 0 56896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1666464484
transform -1 0 50288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1666464484
transform 1 0 1680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1666464484
transform -1 0 57344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1666464484
transform -1 0 1904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1666464484
transform -1 0 34832 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1666464484
transform -1 0 46256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1666464484
transform -1 0 1904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1666464484
transform -1 0 23408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1666464484
transform -1 0 1904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1666464484
transform -1 0 57344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1666464484
transform -1 0 57344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1666464484
transform -1 0 1904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1666464484
transform -1 0 57344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1666464484
transform -1 0 19376 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1666464484
transform -1 0 37520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1666464484
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1666464484
transform -1 0 1904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1666464484
transform -1 0 20832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1666464484
transform -1 0 55216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1666464484
transform -1 0 57344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1666464484
transform -1 0 29456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1666464484
transform -1 0 52192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1666464484
transform -1 0 41552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1666464484
transform -1 0 1904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1666464484
transform -1 0 1904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1666464484
transform -1 0 58240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1666464484
transform 1 0 16464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1666464484
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1666464484
transform -1 0 56448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1666464484
transform 1 0 3248 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1666464484
transform 1 0 34720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1666464484
transform -1 0 4144 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1666464484
transform -1 0 56112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1666464484
transform -1 0 22736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output45_I
timestamp 1666464484
transform -1 0 56448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output46_I
timestamp 1666464484
transform 1 0 56224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1666464484
transform 1 0 3472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1666464484
transform 1 0 3472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1666464484
transform -1 0 20720 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1666464484
transform -1 0 28672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1666464484
transform 1 0 3472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1666464484
transform -1 0 3696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1666464484
transform 1 0 3472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1666464484
transform -1 0 25424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1666464484
transform -1 0 40432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1666464484
transform 1 0 55776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output57_I
timestamp 1666464484
transform -1 0 12880 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output58_I
timestamp 1666464484
transform 1 0 11088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output59_I
timestamp 1666464484
transform 1 0 4368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output60_I
timestamp 1666464484
transform 1 0 56224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1666464484
transform -1 0 3696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1666464484
transform -1 0 16912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output63_I
timestamp 1666464484
transform 1 0 3472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1666464484
transform 1 0 56224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1666464484
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output66_I
timestamp 1666464484
transform 1 0 3472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output67_I
timestamp 1666464484
transform -1 0 49616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1666464484
transform -1 0 7616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 2464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 2688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31
timestamp 1666464484
transform 1 0 4816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1666464484
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1666464484
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 6272 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60
timestamp 1666464484
transform 1 0 8064 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1666464484
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1666464484
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87
timestamp 1666464484
transform 1 0 11088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95
timestamp 1666464484
transform 1 0 11984 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103
timestamp 1666464484
transform 1 0 12880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1666464484
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115
timestamp 1666464484
transform 1 0 14224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119
timestamp 1666464484
transform 1 0 14672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135
timestamp 1666464484
transform 1 0 16464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1666464484
transform 1 0 17472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_159
timestamp 1666464484
transform 1 0 19152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_167
timestamp 1666464484
transform 1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_171
timestamp 1666464484
transform 1 0 20496 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_184
timestamp 1666464484
transform 1 0 21952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_192
timestamp 1666464484
transform 1 0 22848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_194
timestamp 1666464484
transform 1 0 23072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 23408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_205
timestamp 1666464484
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_228
timestamp 1666464484
transform 1 0 26880 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_233
timestamp 1666464484
transform 1 0 27440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_241
timestamp 1666464484
transform 1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_251
timestamp 1666464484
transform 1 0 29456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_259
timestamp 1666464484
transform 1 0 30352 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_275
timestamp 1666464484
transform 1 0 32144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1666464484
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_297
timestamp 1666464484
transform 1 0 34608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_299
timestamp 1666464484
transform 1 0 34832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_356
timestamp 1666464484
transform 1 0 41216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1666464484
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_367
timestamp 1666464484
transform 1 0 42448 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_375
timestamp 1666464484
transform 1 0 43344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_379
timestamp 1666464484
transform 1 0 43792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_381
timestamp 1666464484
transform 1 0 44016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_402
timestamp 1666464484
transform 1 0 46368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_410
timestamp 1666464484
transform 1 0 47264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_414
timestamp 1666464484
transform 1 0 47712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_416
timestamp 1666464484
transform 1 0 47936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1666464484
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_429
timestamp 1666464484
transform 1 0 49392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_433
timestamp 1666464484
transform 1 0 49840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_437
timestamp 1666464484
transform 1 0 50288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_445
timestamp 1666464484
transform 1 0 51184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1666464484
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_457
timestamp 1666464484
transform 1 0 52528 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_473
timestamp 1666464484
transform 1 0 54320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_481
timestamp 1666464484
transform 1 0 55216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_485
timestamp 1666464484
transform 1 0 55664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1666464484
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1666464484
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1666464484
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_17
timestamp 1666464484
transform 1 0 3248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_21
timestamp 1666464484
transform 1 0 3696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_25
timestamp 1666464484
transform 1 0 4144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_29
timestamp 1666464484
transform 1 0 4592 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_61
timestamp 1666464484
transform 1 0 8176 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1666464484
transform 1 0 9072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_81
timestamp 1666464484
transform 1 0 10416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_85
timestamp 1666464484
transform 1 0 10864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_89
timestamp 1666464484
transform 1 0 11312 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_121
timestamp 1666464484
transform 1 0 14896 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_129
timestamp 1666464484
transform 1 0 15792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_133
timestamp 1666464484
transform 1 0 16240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1666464484
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1666464484
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_294
timestamp 1666464484
transform 1 0 34272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_300
timestamp 1666464484
transform 1 0 34944 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_332
timestamp 1666464484
transform 1 0 38528 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_348
timestamp 1666464484
transform 1 0 40320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1666464484
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1666464484
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1666464484
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1666464484
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_492
timestamp 1666464484
transform 1 0 56448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1666464484
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_499
timestamp 1666464484
transform 1 0 57232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_501
timestamp 1666464484
transform 1 0 57456 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_508
timestamp 1666464484
transform 1 0 58240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_17
timestamp 1666464484
transform 1 0 3248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_21
timestamp 1666464484
transform 1 0 3696 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_29
timestamp 1666464484
transform 1 0 4592 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1666464484
transform 1 0 5040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1666464484
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1666464484
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1666464484
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1666464484
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1666464484
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1666464484
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1666464484
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1666464484
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1666464484
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_463
timestamp 1666464484
transform 1 0 53200 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_495
timestamp 1666464484
transform 1 0 56784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_497
timestamp 1666464484
transform 1 0 57008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_500
timestamp 1666464484
transform 1 0 57344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_508
timestamp 1666464484
transform 1 0 58240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_17
timestamp 1666464484
transform 1 0 3248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_21
timestamp 1666464484
transform 1 0 3696 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_53
timestamp 1666464484
transform 1 0 7280 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1666464484
transform 1 0 9072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1666464484
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1666464484
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1666464484
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1666464484
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1666464484
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1666464484
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1666464484
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1666464484
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1666464484
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_499
timestamp 1666464484
transform 1 0 57232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_503
timestamp 1666464484
transform 1 0 57680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_508
timestamp 1666464484
transform 1 0 58240 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1666464484
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1666464484
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1666464484
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1666464484
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1666464484
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1666464484
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1666464484
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1666464484
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_463
timestamp 1666464484
transform 1 0 53200 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_495
timestamp 1666464484
transform 1 0 56784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_503
timestamp 1666464484
transform 1 0 57680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_507
timestamp 1666464484
transform 1 0 58128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1666464484
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1666464484
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1666464484
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1666464484
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1666464484
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1666464484
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1666464484
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1666464484
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1666464484
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_507
timestamp 1666464484
transform 1 0 58128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_5
timestamp 1666464484
transform 1 0 1904 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_21
timestamp 1666464484
transform 1 0 3696 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_29
timestamp 1666464484
transform 1 0 4592 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_33
timestamp 1666464484
transform 1 0 5040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1666464484
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1666464484
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1666464484
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1666464484
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1666464484
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_463
timestamp 1666464484
transform 1 0 53200 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_495
timestamp 1666464484
transform 1 0 56784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_497
timestamp 1666464484
transform 1 0 57008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_500
timestamp 1666464484
transform 1 0 57344 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_508
timestamp 1666464484
transform 1 0 58240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_9
timestamp 1666464484
transform 1 0 2352 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_41
timestamp 1666464484
transform 1 0 5936 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_57
timestamp 1666464484
transform 1 0 7728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_65
timestamp 1666464484
transform 1 0 8624 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1666464484
transform 1 0 9072 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1666464484
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1666464484
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1666464484
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1666464484
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1666464484
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1666464484
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_499
timestamp 1666464484
transform 1 0 57232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_507
timestamp 1666464484
transform 1 0 58128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1666464484
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1666464484
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1666464484
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_463
timestamp 1666464484
transform 1 0 53200 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_495
timestamp 1666464484
transform 1 0 56784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_503
timestamp 1666464484
transform 1 0 57680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_507
timestamp 1666464484
transform 1 0 58128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1666464484
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1666464484
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1666464484
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1666464484
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1666464484
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1666464484
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1666464484
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1666464484
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1666464484
transform 1 0 57232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_507
timestamp 1666464484
transform 1 0 58128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1666464484
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1666464484
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1666464484
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1666464484
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1666464484
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_463
timestamp 1666464484
transform 1 0 53200 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_479
timestamp 1666464484
transform 1 0 54992 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_487
timestamp 1666464484
transform 1 0 55888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_489
timestamp 1666464484
transform 1 0 56112 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_492
timestamp 1666464484
transform 1 0 56448 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_508
timestamp 1666464484
transform 1 0 58240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_17
timestamp 1666464484
transform 1 0 3248 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_21
timestamp 1666464484
transform 1 0 3696 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_53
timestamp 1666464484
transform 1 0 7280 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1666464484
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1666464484
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1666464484
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1666464484
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1666464484
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1666464484
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_499
timestamp 1666464484
transform 1 0 57232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_507
timestamp 1666464484
transform 1 0 58128 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1666464484
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_463
timestamp 1666464484
transform 1 0 53200 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_495
timestamp 1666464484
transform 1 0 56784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_503
timestamp 1666464484
transform 1 0 57680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_507
timestamp 1666464484
transform 1 0 58128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1666464484
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1666464484
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1666464484
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1666464484
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1666464484
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_499
timestamp 1666464484
transform 1 0 57232 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_507
timestamp 1666464484
transform 1 0 58128 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_5
timestamp 1666464484
transform 1 0 1904 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_21
timestamp 1666464484
transform 1 0 3696 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_29
timestamp 1666464484
transform 1 0 4592 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1666464484
transform 1 0 5040 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1666464484
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1666464484
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_463
timestamp 1666464484
transform 1 0 53200 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_479
timestamp 1666464484
transform 1 0 54992 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_487
timestamp 1666464484
transform 1 0 55888 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_489
timestamp 1666464484
transform 1 0 56112 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_492
timestamp 1666464484
transform 1 0 56448 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_508
timestamp 1666464484
transform 1 0 58240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_9
timestamp 1666464484
transform 1 0 2352 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_41
timestamp 1666464484
transform 1 0 5936 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_57
timestamp 1666464484
transform 1 0 7728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_65
timestamp 1666464484
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1666464484
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1666464484
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1666464484
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1666464484
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1666464484
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1666464484
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_499
timestamp 1666464484
transform 1 0 57232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_507
timestamp 1666464484
transform 1 0 58128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1666464484
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1666464484
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1666464484
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_463
timestamp 1666464484
transform 1 0 53200 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_495
timestamp 1666464484
transform 1 0 56784 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_503
timestamp 1666464484
transform 1 0 57680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_507
timestamp 1666464484
transform 1 0 58128 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_5
timestamp 1666464484
transform 1 0 1904 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_69
timestamp 1666464484
transform 1 0 9072 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1666464484
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1666464484
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1666464484
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1666464484
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1666464484
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1666464484
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_499
timestamp 1666464484
transform 1 0 57232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_507
timestamp 1666464484
transform 1 0 58128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_9
timestamp 1666464484
transform 1 0 2352 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_25
timestamp 1666464484
transform 1 0 4144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1666464484
transform 1 0 5040 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1666464484
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1666464484
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_463
timestamp 1666464484
transform 1 0 53200 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_495
timestamp 1666464484
transform 1 0 56784 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_497
timestamp 1666464484
transform 1 0 57008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_500
timestamp 1666464484
transform 1 0 57344 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_508
timestamp 1666464484
transform 1 0 58240 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1666464484
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1666464484
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1666464484
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1666464484
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_499
timestamp 1666464484
transform 1 0 57232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_507
timestamp 1666464484
transform 1 0 58128 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1666464484
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1666464484
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_463
timestamp 1666464484
transform 1 0 53200 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_495
timestamp 1666464484
transform 1 0 56784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_503
timestamp 1666464484
transform 1 0 57680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_507
timestamp 1666464484
transform 1 0 58128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1666464484
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1666464484
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1666464484
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1666464484
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1666464484
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_499
timestamp 1666464484
transform 1 0 57232 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_507
timestamp 1666464484
transform 1 0 58128 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_18
timestamp 1666464484
transform 1 0 3360 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_28
timestamp 1666464484
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_32
timestamp 1666464484
transform 1 0 4928 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1666464484
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1666464484
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_463
timestamp 1666464484
transform 1 0 53200 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_495
timestamp 1666464484
transform 1 0 56784 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_497
timestamp 1666464484
transform 1 0 57008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_500
timestamp 1666464484
transform 1 0 57344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_508
timestamp 1666464484
transform 1 0 58240 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_17
timestamp 1666464484
transform 1 0 3248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_21
timestamp 1666464484
transform 1 0 3696 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_53
timestamp 1666464484
transform 1 0 7280 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_69
timestamp 1666464484
transform 1 0 9072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_91
timestamp 1666464484
transform 1 0 11536 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_123
timestamp 1666464484
transform 1 0 15120 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_139
timestamp 1666464484
transform 1 0 16912 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1666464484
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1666464484
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1666464484
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1666464484
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1666464484
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_499
timestamp 1666464484
transform 1 0 57232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_507
timestamp 1666464484
transform 1 0 58128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1666464484
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_69
timestamp 1666464484
transform 1 0 9072 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_71
timestamp 1666464484
transform 1 0 9296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_74
timestamp 1666464484
transform 1 0 9632 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_89
timestamp 1666464484
transform 1 0 11312 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_95
timestamp 1666464484
transform 1 0 11984 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_99
timestamp 1666464484
transform 1 0 12432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_103
timestamp 1666464484
transform 1 0 12880 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1666464484
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1666464484
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_463
timestamp 1666464484
transform 1 0 53200 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_495
timestamp 1666464484
transform 1 0 56784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_503
timestamp 1666464484
transform 1 0 57680 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_505
timestamp 1666464484
transform 1 0 57904 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_508
timestamp 1666464484
transform 1 0 58240 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_86
timestamp 1666464484
transform 1 0 10976 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_90
timestamp 1666464484
transform 1 0 11424 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_94
timestamp 1666464484
transform 1 0 11872 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_126
timestamp 1666464484
transform 1 0 15456 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_134
timestamp 1666464484
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_138
timestamp 1666464484
transform 1 0 16800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_153
timestamp 1666464484
transform 1 0 18480 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_157
timestamp 1666464484
transform 1 0 18928 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_161
timestamp 1666464484
transform 1 0 19376 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_179
timestamp 1666464484
transform 1 0 21392 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_183
timestamp 1666464484
transform 1 0 21840 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_196
timestamp 1666464484
transform 1 0 23296 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_200
timestamp 1666464484
transform 1 0 23744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1666464484
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1666464484
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1666464484
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_499
timestamp 1666464484
transform 1 0 57232 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_501
timestamp 1666464484
transform 1 0 57456 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_508
timestamp 1666464484
transform 1 0 58240 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_17
timestamp 1666464484
transform 1 0 3248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_21
timestamp 1666464484
transform 1 0 3696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_29
timestamp 1666464484
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_33
timestamp 1666464484
transform 1 0 5040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_148
timestamp 1666464484
transform 1 0 17920 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_152
timestamp 1666464484
transform 1 0 18368 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_156
timestamp 1666464484
transform 1 0 18816 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_183
timestamp 1666464484
transform 1 0 21840 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_187
timestamp 1666464484
transform 1 0 22288 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_221
timestamp 1666464484
transform 1 0 26096 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_225
timestamp 1666464484
transform 1 0 26544 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_241
timestamp 1666464484
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_245
timestamp 1666464484
transform 1 0 28784 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1666464484
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1666464484
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_463
timestamp 1666464484
transform 1 0 53200 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_495
timestamp 1666464484
transform 1 0 56784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_503
timestamp 1666464484
transform 1 0 57680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_507
timestamp 1666464484
transform 1 0 58128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_77
timestamp 1666464484
transform 1 0 9968 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_81
timestamp 1666464484
transform 1 0 10416 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_83
timestamp 1666464484
transform 1 0 10640 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_91
timestamp 1666464484
transform 1 0 11536 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_95
timestamp 1666464484
transform 1 0 11984 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_99
timestamp 1666464484
transform 1 0 12432 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_131
timestamp 1666464484
transform 1 0 16016 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_139
timestamp 1666464484
transform 1 0 16912 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_160
timestamp 1666464484
transform 1 0 19264 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_166
timestamp 1666464484
transform 1 0 19936 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_184
timestamp 1666464484
transform 1 0 21952 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_190
timestamp 1666464484
transform 1 0 22624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_194
timestamp 1666464484
transform 1 0 23072 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_197
timestamp 1666464484
transform 1 0 23408 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_201
timestamp 1666464484
transform 1 0 23856 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_210
timestamp 1666464484
transform 1 0 24864 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_223
timestamp 1666464484
transform 1 0 26320 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_227
timestamp 1666464484
transform 1 0 26768 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_230
timestamp 1666464484
transform 1 0 27104 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_234
timestamp 1666464484
transform 1 0 27552 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_238
timestamp 1666464484
transform 1 0 28000 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_247
timestamp 1666464484
transform 1 0 29008 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1666464484
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1666464484
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1666464484
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1666464484
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1666464484
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_499
timestamp 1666464484
transform 1 0 57232 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_507
timestamp 1666464484
transform 1 0 58128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1666464484
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_69
timestamp 1666464484
transform 1 0 9072 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_79
timestamp 1666464484
transform 1 0 10192 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_93
timestamp 1666464484
transform 1 0 11760 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_191
timestamp 1666464484
transform 1 0 22736 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_195
timestamp 1666464484
transform 1 0 23184 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_199
timestamp 1666464484
transform 1 0 23632 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_206
timestamp 1666464484
transform 1 0 24416 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_210
timestamp 1666464484
transform 1 0 24864 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_242
timestamp 1666464484
transform 1 0 28448 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_246
timestamp 1666464484
transform 1 0 28896 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1666464484
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1666464484
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_463
timestamp 1666464484
transform 1 0 53200 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_479
timestamp 1666464484
transform 1 0 54992 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_487
timestamp 1666464484
transform 1 0 55888 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_489
timestamp 1666464484
transform 1 0 56112 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_492
timestamp 1666464484
transform 1 0 56448 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_508
timestamp 1666464484
transform 1 0 58240 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_77
timestamp 1666464484
transform 1 0 9968 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_81
timestamp 1666464484
transform 1 0 10416 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_91
timestamp 1666464484
transform 1 0 11536 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_97
timestamp 1666464484
transform 1 0 12208 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_101
timestamp 1666464484
transform 1 0 12656 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_133
timestamp 1666464484
transform 1 0 16240 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_176
timestamp 1666464484
transform 1 0 21056 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_192
timestamp 1666464484
transform 1 0 22848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_196
timestamp 1666464484
transform 1 0 23296 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_200
timestamp 1666464484
transform 1 0 23744 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_204
timestamp 1666464484
transform 1 0 24192 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_218
timestamp 1666464484
transform 1 0 25760 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_226
timestamp 1666464484
transform 1 0 26656 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_234
timestamp 1666464484
transform 1 0 27552 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_238
timestamp 1666464484
transform 1 0 28000 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_270
timestamp 1666464484
transform 1 0 31584 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_274
timestamp 1666464484
transform 1 0 32032 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_277
timestamp 1666464484
transform 1 0 32368 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 32816 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_366
timestamp 1666464484
transform 1 0 42336 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_370
timestamp 1666464484
transform 1 0 42784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_374
timestamp 1666464484
transform 1 0 43232 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_406
timestamp 1666464484
transform 1 0 46816 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_422
timestamp 1666464484
transform 1 0 48608 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1666464484
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1666464484
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1666464484
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_499
timestamp 1666464484
transform 1 0 57232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_507
timestamp 1666464484
transform 1 0 58128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_17
timestamp 1666464484
transform 1 0 3248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_21
timestamp 1666464484
transform 1 0 3696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_29
timestamp 1666464484
transform 1 0 4592 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_33
timestamp 1666464484
transform 1 0 5040 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_69
timestamp 1666464484
transform 1 0 9072 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_85
timestamp 1666464484
transform 1 0 10864 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_87
timestamp 1666464484
transform 1 0 11088 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_94
timestamp 1666464484
transform 1 0 11872 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_98
timestamp 1666464484
transform 1 0 12320 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_140
timestamp 1666464484
transform 1 0 17024 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_142
timestamp 1666464484
transform 1 0 17248 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_145
timestamp 1666464484
transform 1 0 17584 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_149
timestamp 1666464484
transform 1 0 18032 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_153
timestamp 1666464484
transform 1 0 18480 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_166
timestamp 1666464484
transform 1 0 19936 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_170
timestamp 1666464484
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_174
timestamp 1666464484
transform 1 0 20832 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_187
timestamp 1666464484
transform 1 0 22288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_191
timestamp 1666464484
transform 1 0 22736 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_200
timestamp 1666464484
transform 1 0 23744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_216
timestamp 1666464484
transform 1 0 25536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_222
timestamp 1666464484
transform 1 0 26208 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_226
timestamp 1666464484
transform 1 0 26656 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_246
timestamp 1666464484
transform 1 0 28896 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_253
timestamp 1666464484
transform 1 0 29680 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_261
timestamp 1666464484
transform 1 0 30576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_265
timestamp 1666464484
transform 1 0 31024 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_269
timestamp 1666464484
transform 1 0 31472 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_273
timestamp 1666464484
transform 1 0 31920 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_293
timestamp 1666464484
transform 1 0 34160 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_309
timestamp 1666464484
transform 1 0 35952 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_317
timestamp 1666464484
transform 1 0 36848 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1666464484
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1666464484
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_463
timestamp 1666464484
transform 1 0 53200 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_495
timestamp 1666464484
transform 1 0 56784 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_503
timestamp 1666464484
transform 1 0 57680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_507
timestamp 1666464484
transform 1 0 58128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_34
timestamp 1666464484
transform 1 0 5152 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_38
timestamp 1666464484
transform 1 0 5600 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_46
timestamp 1666464484
transform 1 0 6496 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_50
timestamp 1666464484
transform 1 0 6944 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_54
timestamp 1666464484
transform 1 0 7392 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1666464484
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_89
timestamp 1666464484
transform 1 0 11312 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_93
timestamp 1666464484
transform 1 0 11760 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_97
timestamp 1666464484
transform 1 0 12208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_101
timestamp 1666464484
transform 1 0 12656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_104
timestamp 1666464484
transform 1 0 12992 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_136
timestamp 1666464484
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_140
timestamp 1666464484
transform 1 0 17024 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_147
timestamp 1666464484
transform 1 0 17808 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_179
timestamp 1666464484
transform 1 0 21392 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_187
timestamp 1666464484
transform 1 0 22288 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_191
timestamp 1666464484
transform 1 0 22736 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_193
timestamp 1666464484
transform 1 0 22960 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_202
timestamp 1666464484
transform 1 0 23968 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_206
timestamp 1666464484
transform 1 0 24416 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_210
timestamp 1666464484
transform 1 0 24864 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_231
timestamp 1666464484
transform 1 0 27216 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_239
timestamp 1666464484
transform 1 0 28112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_241
timestamp 1666464484
transform 1 0 28336 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_247
timestamp 1666464484
transform 1 0 29008 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_251
timestamp 1666464484
transform 1 0 29456 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1666464484
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1666464484
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1666464484
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1666464484
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1666464484
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_499
timestamp 1666464484
transform 1 0 57232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_507
timestamp 1666464484
transform 1 0 58128 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1666464484
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_69
timestamp 1666464484
transform 1 0 9072 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_85
timestamp 1666464484
transform 1 0 10864 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_91
timestamp 1666464484
transform 1 0 11536 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_93
timestamp 1666464484
transform 1 0 11760 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_102
timestamp 1666464484
transform 1 0 12768 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_111
timestamp 1666464484
transform 1 0 13776 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_127
timestamp 1666464484
transform 1 0 15568 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_131
timestamp 1666464484
transform 1 0 16016 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_141
timestamp 1666464484
transform 1 0 17136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_145
timestamp 1666464484
transform 1 0 17584 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_148
timestamp 1666464484
transform 1 0 17920 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_159
timestamp 1666464484
transform 1 0 19152 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_163
timestamp 1666464484
transform 1 0 19600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_171
timestamp 1666464484
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_175
timestamp 1666464484
transform 1 0 20944 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_187
timestamp 1666464484
transform 1 0 22288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_202
timestamp 1666464484
transform 1 0 23968 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_206
timestamp 1666464484
transform 1 0 24416 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_210
timestamp 1666464484
transform 1 0 24864 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_218
timestamp 1666464484
transform 1 0 25760 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_222
timestamp 1666464484
transform 1 0 26208 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_226
timestamp 1666464484
transform 1 0 26656 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_240
timestamp 1666464484
transform 1 0 28224 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_244
timestamp 1666464484
transform 1 0 28672 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_282
timestamp 1666464484
transform 1 0 32928 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_284
timestamp 1666464484
transform 1 0 33152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_287
timestamp 1666464484
transform 1 0 33488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_291
timestamp 1666464484
transform 1 0 33936 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_295
timestamp 1666464484
transform 1 0 34384 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_299
timestamp 1666464484
transform 1 0 34832 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_311
timestamp 1666464484
transform 1 0 36176 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_325
timestamp 1666464484
transform 1 0 37744 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_327
timestamp 1666464484
transform 1 0 37968 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_330
timestamp 1666464484
transform 1 0 38304 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_334
timestamp 1666464484
transform 1 0 38752 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_346
timestamp 1666464484
transform 1 0 40096 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_350
timestamp 1666464484
transform 1 0 40544 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_354
timestamp 1666464484
transform 1 0 40992 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_362
timestamp 1666464484
transform 1 0 41888 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_366
timestamp 1666464484
transform 1 0 42336 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_382
timestamp 1666464484
transform 1 0 44128 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1666464484
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_463
timestamp 1666464484
transform 1 0 53200 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_495
timestamp 1666464484
transform 1 0 56784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_503
timestamp 1666464484
transform 1 0 57680 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_505
timestamp 1666464484
transform 1 0 57904 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_508
timestamp 1666464484
transform 1 0 58240 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_5
timestamp 1666464484
transform 1 0 1904 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_37
timestamp 1666464484
transform 1 0 5488 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_53
timestamp 1666464484
transform 1 0 7280 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_61
timestamp 1666464484
transform 1 0 8176 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_65
timestamp 1666464484
transform 1 0 8624 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1666464484
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_89
timestamp 1666464484
transform 1 0 11312 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_99
timestamp 1666464484
transform 1 0 12432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_107
timestamp 1666464484
transform 1 0 13328 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_111
timestamp 1666464484
transform 1 0 13776 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_113
timestamp 1666464484
transform 1 0 14000 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_116
timestamp 1666464484
transform 1 0 14336 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_132
timestamp 1666464484
transform 1 0 16128 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_136
timestamp 1666464484
transform 1 0 16576 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_138
timestamp 1666464484
transform 1 0 16800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_147
timestamp 1666464484
transform 1 0 17808 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_160
timestamp 1666464484
transform 1 0 19264 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_164
timestamp 1666464484
transform 1 0 19712 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_168
timestamp 1666464484
transform 1 0 20160 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_172
timestamp 1666464484
transform 1 0 20608 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_180
timestamp 1666464484
transform 1 0 21504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_184
timestamp 1666464484
transform 1 0 21952 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_188
timestamp 1666464484
transform 1 0 22400 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_198
timestamp 1666464484
transform 1 0 23520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_202
timestamp 1666464484
transform 1 0 23968 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_206
timestamp 1666464484
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_224
timestamp 1666464484
transform 1 0 26432 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_256
timestamp 1666464484
transform 1 0 30016 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_272
timestamp 1666464484
transform 1 0 31808 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_274
timestamp 1666464484
transform 1 0 32032 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_277
timestamp 1666464484
transform 1 0 32368 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_293
timestamp 1666464484
transform 1 0 34160 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_297
timestamp 1666464484
transform 1 0 34608 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_329
timestamp 1666464484
transform 1 0 38192 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_345
timestamp 1666464484
transform 1 0 39984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_353
timestamp 1666464484
transform 1 0 40880 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1666464484
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1666464484
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1666464484
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1666464484
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1666464484
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_499
timestamp 1666464484
transform 1 0 57232 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_501
timestamp 1666464484
transform 1 0 57456 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_508
timestamp 1666464484
transform 1 0 58240 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_9
timestamp 1666464484
transform 1 0 2352 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_25
timestamp 1666464484
transform 1 0 4144 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_33
timestamp 1666464484
transform 1 0 5040 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_44
timestamp 1666464484
transform 1 0 6272 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_48
timestamp 1666464484
transform 1 0 6720 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_56
timestamp 1666464484
transform 1 0 7616 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_59
timestamp 1666464484
transform 1 0 7952 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_67
timestamp 1666464484
transform 1 0 8848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_81
timestamp 1666464484
transform 1 0 10416 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_85
timestamp 1666464484
transform 1 0 10864 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_91
timestamp 1666464484
transform 1 0 11536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_95
timestamp 1666464484
transform 1 0 11984 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_100
timestamp 1666464484
transform 1 0 12544 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_104
timestamp 1666464484
transform 1 0 12992 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_114
timestamp 1666464484
transform 1 0 14112 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_118
timestamp 1666464484
transform 1 0 14560 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_120
timestamp 1666464484
transform 1 0 14784 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_123
timestamp 1666464484
transform 1 0 15120 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_133
timestamp 1666464484
transform 1 0 16240 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_139
timestamp 1666464484
transform 1 0 16912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_143
timestamp 1666464484
transform 1 0 17360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_157
timestamp 1666464484
transform 1 0 18928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_170
timestamp 1666464484
transform 1 0 20384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_182
timestamp 1666464484
transform 1 0 21728 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1666464484
transform 1 0 28896 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_268
timestamp 1666464484
transform 1 0 31360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_272
timestamp 1666464484
transform 1 0 31808 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_281
timestamp 1666464484
transform 1 0 32816 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_313
timestamp 1666464484
transform 1 0 36400 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1666464484
transform 1 0 36848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1666464484
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1666464484
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_463
timestamp 1666464484
transform 1 0 53200 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_495
timestamp 1666464484
transform 1 0 56784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_503
timestamp 1666464484
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_507
timestamp 1666464484
transform 1 0 58128 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_18
timestamp 1666464484
transform 1 0 3360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_26
timestamp 1666464484
transform 1 0 4256 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_28
timestamp 1666464484
transform 1 0 4480 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_31
timestamp 1666464484
transform 1 0 4816 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_39
timestamp 1666464484
transform 1 0 5712 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_43
timestamp 1666464484
transform 1 0 6160 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_59
timestamp 1666464484
transform 1 0 7952 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_67
timestamp 1666464484
transform 1 0 8848 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_83
timestamp 1666464484
transform 1 0 10640 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_87
timestamp 1666464484
transform 1 0 11088 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_91
timestamp 1666464484
transform 1 0 11536 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_98
timestamp 1666464484
transform 1 0 12320 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_112
timestamp 1666464484
transform 1 0 13888 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_128
timestamp 1666464484
transform 1 0 15680 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_136
timestamp 1666464484
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_140
timestamp 1666464484
transform 1 0 17024 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_152
timestamp 1666464484
transform 1 0 18368 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_156
timestamp 1666464484
transform 1 0 18816 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_159
timestamp 1666464484
transform 1 0 19152 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_191
timestamp 1666464484
transform 1 0 22736 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_207
timestamp 1666464484
transform 1 0 24528 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_211
timestamp 1666464484
transform 1 0 24976 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_231
timestamp 1666464484
transform 1 0 27216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_235
timestamp 1666464484
transform 1 0 27664 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_237
timestamp 1666464484
transform 1 0 27888 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_240
timestamp 1666464484
transform 1 0 28224 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_248
timestamp 1666464484
transform 1 0 29120 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_252
timestamp 1666464484
transform 1 0 29568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_318
timestamp 1666464484
transform 1 0 36960 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_324
timestamp 1666464484
transform 1 0 37632 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_340
timestamp 1666464484
transform 1 0 39424 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_348
timestamp 1666464484
transform 1 0 40320 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_352
timestamp 1666464484
transform 1 0 40768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_360
timestamp 1666464484
transform 1 0 41664 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_424
timestamp 1666464484
transform 1 0 48832 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1666464484
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1666464484
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1666464484
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_499
timestamp 1666464484
transform 1 0 57232 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_507
timestamp 1666464484
transform 1 0 58128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_69
timestamp 1666464484
transform 1 0 9072 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_85
timestamp 1666464484
transform 1 0 10864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_88
timestamp 1666464484
transform 1 0 11200 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_96
timestamp 1666464484
transform 1 0 12096 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_100
timestamp 1666464484
transform 1 0 12544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_104
timestamp 1666464484
transform 1 0 12992 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_124
timestamp 1666464484
transform 1 0 15232 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_128
timestamp 1666464484
transform 1 0 15680 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_130
timestamp 1666464484
transform 1 0 15904 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_133
timestamp 1666464484
transform 1 0 16240 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_142
timestamp 1666464484
transform 1 0 17248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_146
timestamp 1666464484
transform 1 0 17696 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_150
timestamp 1666464484
transform 1 0 18144 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_166
timestamp 1666464484
transform 1 0 19936 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_174
timestamp 1666464484
transform 1 0 20832 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_183
timestamp 1666464484
transform 1 0 21840 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_186
timestamp 1666464484
transform 1 0 22176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 23072 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_196
timestamp 1666464484
transform 1 0 23296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_203
timestamp 1666464484
transform 1 0 24080 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_207
timestamp 1666464484
transform 1 0 24528 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_211
timestamp 1666464484
transform 1 0 24976 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_229
timestamp 1666464484
transform 1 0 26992 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_233
timestamp 1666464484
transform 1 0 27440 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_241
timestamp 1666464484
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_245
timestamp 1666464484
transform 1 0 28784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_258
timestamp 1666464484
transform 1 0 30240 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_265
timestamp 1666464484
transform 1 0 31024 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_269
timestamp 1666464484
transform 1 0 31472 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_273
timestamp 1666464484
transform 1 0 31920 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_289
timestamp 1666464484
transform 1 0 33712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_291
timestamp 1666464484
transform 1 0 33936 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_294
timestamp 1666464484
transform 1 0 34272 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_302
timestamp 1666464484
transform 1 0 35168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_308
timestamp 1666464484
transform 1 0 35840 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_323
timestamp 1666464484
transform 1 0 37520 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_334
timestamp 1666464484
transform 1 0 38752 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_342
timestamp 1666464484
transform 1 0 39648 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_346
timestamp 1666464484
transform 1 0 40096 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_350
timestamp 1666464484
transform 1 0 40544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_354
timestamp 1666464484
transform 1 0 40992 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_359
timestamp 1666464484
transform 1 0 41552 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_363
timestamp 1666464484
transform 1 0 42000 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_379
timestamp 1666464484
transform 1 0 43792 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_387
timestamp 1666464484
transform 1 0 44688 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1666464484
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_463
timestamp 1666464484
transform 1 0 53200 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_495
timestamp 1666464484
transform 1 0 56784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_503
timestamp 1666464484
transform 1 0 57680 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_508
timestamp 1666464484
transform 1 0 58240 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_17
timestamp 1666464484
transform 1 0 3248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_21
timestamp 1666464484
transform 1 0 3696 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_53
timestamp 1666464484
transform 1 0 7280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_69
timestamp 1666464484
transform 1 0 9072 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_86
timestamp 1666464484
transform 1 0 10976 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_93
timestamp 1666464484
transform 1 0 11760 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_103
timestamp 1666464484
transform 1 0 12880 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_107
timestamp 1666464484
transform 1 0 13328 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_139
timestamp 1666464484
transform 1 0 16912 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_176
timestamp 1666464484
transform 1 0 21056 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_178
timestamp 1666464484
transform 1 0 21280 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_184
timestamp 1666464484
transform 1 0 21952 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_194
timestamp 1666464484
transform 1 0 23072 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_198
timestamp 1666464484
transform 1 0 23520 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_202
timestamp 1666464484
transform 1 0 23968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_227
timestamp 1666464484
transform 1 0 26768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_241
timestamp 1666464484
transform 1 0 28336 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_245
timestamp 1666464484
transform 1 0 28784 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_277
timestamp 1666464484
transform 1 0 32368 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_281
timestamp 1666464484
transform 1 0 32816 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_292
timestamp 1666464484
transform 1 0 34048 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_299
timestamp 1666464484
transform 1 0 34832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_306
timestamp 1666464484
transform 1 0 35616 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_310
timestamp 1666464484
transform 1 0 36064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_314
timestamp 1666464484
transform 1 0 36512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_318
timestamp 1666464484
transform 1 0 36960 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_323
timestamp 1666464484
transform 1 0 37520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_333
timestamp 1666464484
transform 1 0 38640 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 39088 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_339
timestamp 1666464484
transform 1 0 39312 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_348
timestamp 1666464484
transform 1 0 40320 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_352
timestamp 1666464484
transform 1 0 40768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_361
timestamp 1666464484
transform 1 0 41776 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_371
timestamp 1666464484
transform 1 0 42896 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_403
timestamp 1666464484
transform 1 0 46480 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_419
timestamp 1666464484
transform 1 0 48272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_423
timestamp 1666464484
transform 1 0 48720 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1666464484
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1666464484
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1666464484
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1666464484
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_499
timestamp 1666464484
transform 1 0 57232 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_507
timestamp 1666464484
transform 1 0 58128 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_69
timestamp 1666464484
transform 1 0 9072 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_85
timestamp 1666464484
transform 1 0 10864 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_89
timestamp 1666464484
transform 1 0 11312 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_92
timestamp 1666464484
transform 1 0 11648 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_96
timestamp 1666464484
transform 1 0 12096 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_104
timestamp 1666464484
transform 1 0 12992 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_124
timestamp 1666464484
transform 1 0 15232 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_134
timestamp 1666464484
transform 1 0 16352 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_144
timestamp 1666464484
transform 1 0 17472 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_195
timestamp 1666464484
transform 1 0 23184 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_199
timestamp 1666464484
transform 1 0 23632 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_201
timestamp 1666464484
transform 1 0 23856 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_204
timestamp 1666464484
transform 1 0 24192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_208
timestamp 1666464484
transform 1 0 24640 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_212
timestamp 1666464484
transform 1 0 25088 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_225
timestamp 1666464484
transform 1 0 26544 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_232
timestamp 1666464484
transform 1 0 27328 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_238
timestamp 1666464484
transform 1 0 28000 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_242
timestamp 1666464484
transform 1 0 28448 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_244
timestamp 1666464484
transform 1 0 28672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_256
timestamp 1666464484
transform 1 0 30016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_260
timestamp 1666464484
transform 1 0 30464 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_268
timestamp 1666464484
transform 1 0 31360 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_270
timestamp 1666464484
transform 1 0 31584 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_273
timestamp 1666464484
transform 1 0 31920 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_281
timestamp 1666464484
transform 1 0 32816 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_285
timestamp 1666464484
transform 1 0 33264 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_289
timestamp 1666464484
transform 1 0 33712 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_291
timestamp 1666464484
transform 1 0 33936 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_306
timestamp 1666464484
transform 1 0 35616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_334
timestamp 1666464484
transform 1 0 38752 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_338
timestamp 1666464484
transform 1 0 39200 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_348
timestamp 1666464484
transform 1 0 40320 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_356
timestamp 1666464484
transform 1 0 41216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_360
timestamp 1666464484
transform 1 0 41664 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_365
timestamp 1666464484
transform 1 0 42224 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_369
timestamp 1666464484
transform 1 0 42672 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_424
timestamp 1666464484
transform 1 0 48832 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_428
timestamp 1666464484
transform 1 0 49280 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_437
timestamp 1666464484
transform 1 0 50288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_441
timestamp 1666464484
transform 1 0 50736 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_457
timestamp 1666464484
transform 1 0 52528 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_463
timestamp 1666464484
transform 1 0 53200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_495
timestamp 1666464484
transform 1 0 56784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_503
timestamp 1666464484
transform 1 0 57680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1666464484
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_18
timestamp 1666464484
transform 1 0 3360 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_26
timestamp 1666464484
transform 1 0 4256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_28
timestamp 1666464484
transform 1 0 4480 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_35
timestamp 1666464484
transform 1 0 5264 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_39
timestamp 1666464484
transform 1 0 5712 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_55
timestamp 1666464484
transform 1 0 7504 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_57
timestamp 1666464484
transform 1 0 7728 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_62
timestamp 1666464484
transform 1 0 8288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_86
timestamp 1666464484
transform 1 0 10976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_90
timestamp 1666464484
transform 1 0 11424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_94
timestamp 1666464484
transform 1 0 11872 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_126
timestamp 1666464484
transform 1 0 15456 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_160
timestamp 1666464484
transform 1 0 19264 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_168
timestamp 1666464484
transform 1 0 20160 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_172
timestamp 1666464484
transform 1 0 20608 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_204
timestamp 1666464484
transform 1 0 24192 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_223
timestamp 1666464484
transform 1 0 26320 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_227
timestamp 1666464484
transform 1 0 26768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_231
timestamp 1666464484
transform 1 0 27216 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_263
timestamp 1666464484
transform 1 0 30800 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_292
timestamp 1666464484
transform 1 0 34048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_302
timestamp 1666464484
transform 1 0 35168 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_308
timestamp 1666464484
transform 1 0 35840 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_312
timestamp 1666464484
transform 1 0 36288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_316
timestamp 1666464484
transform 1 0 36736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_320
timestamp 1666464484
transform 1 0 37184 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_324
timestamp 1666464484
transform 1 0 37632 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_328
timestamp 1666464484
transform 1 0 38080 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_344
timestamp 1666464484
transform 1 0 39872 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_352
timestamp 1666464484
transform 1 0 40768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_389
timestamp 1666464484
transform 1 0 44912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_393
timestamp 1666464484
transform 1 0 45360 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_401
timestamp 1666464484
transform 1 0 46256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_405
timestamp 1666464484
transform 1 0 46704 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1666464484
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1666464484
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1666464484
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1666464484
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1666464484
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_499
timestamp 1666464484
transform 1 0 57232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_507
timestamp 1666464484
transform 1 0 58128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1666464484
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_53
timestamp 1666464484
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_61
timestamp 1666464484
transform 1 0 8176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_65
timestamp 1666464484
transform 1 0 8624 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_67
timestamp 1666464484
transform 1 0 8848 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_70
timestamp 1666464484
transform 1 0 9184 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_76
timestamp 1666464484
transform 1 0 9856 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_86
timestamp 1666464484
transform 1 0 10976 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_90
timestamp 1666464484
transform 1 0 11424 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_99
timestamp 1666464484
transform 1 0 12432 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_103
timestamp 1666464484
transform 1 0 12880 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_116
timestamp 1666464484
transform 1 0 14336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_132
timestamp 1666464484
transform 1 0 16128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_136
timestamp 1666464484
transform 1 0 16576 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_138
timestamp 1666464484
transform 1 0 16800 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 17136 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_155
timestamp 1666464484
transform 1 0 18704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_163
timestamp 1666464484
transform 1 0 19600 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_167
timestamp 1666464484
transform 1 0 20048 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_169
timestamp 1666464484
transform 1 0 20272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_172
timestamp 1666464484
transform 1 0 20608 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_190
timestamp 1666464484
transform 1 0 22624 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 23072 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_198
timestamp 1666464484
transform 1 0 23520 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_202
timestamp 1666464484
transform 1 0 23968 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_206
timestamp 1666464484
transform 1 0 24416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_220
timestamp 1666464484
transform 1 0 25984 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_224
timestamp 1666464484
transform 1 0 26432 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_228
timestamp 1666464484
transform 1 0 26880 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_244
timestamp 1666464484
transform 1 0 28672 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_255
timestamp 1666464484
transform 1 0 29904 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_259
timestamp 1666464484
transform 1 0 30352 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_275
timestamp 1666464484
transform 1 0 32144 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_283
timestamp 1666464484
transform 1 0 33040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_287
timestamp 1666464484
transform 1 0 33488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_295
timestamp 1666464484
transform 1 0 34384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_304
timestamp 1666464484
transform 1 0 35392 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_308
timestamp 1666464484
transform 1 0 35840 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_312
timestamp 1666464484
transform 1 0 36288 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_316
timestamp 1666464484
transform 1 0 36736 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_339
timestamp 1666464484
transform 1 0 39312 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_351
timestamp 1666464484
transform 1 0 40656 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_383
timestamp 1666464484
transform 1 0 44240 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_402
timestamp 1666464484
transform 1 0 46368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_406
timestamp 1666464484
transform 1 0 46816 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_422
timestamp 1666464484
transform 1 0 48608 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_430
timestamp 1666464484
transform 1 0 49504 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_434
timestamp 1666464484
transform 1 0 49952 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_436
timestamp 1666464484
transform 1 0 50176 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_439
timestamp 1666464484
transform 1 0 50512 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_455
timestamp 1666464484
transform 1 0 52304 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_459
timestamp 1666464484
transform 1 0 52752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_463
timestamp 1666464484
transform 1 0 53200 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_479
timestamp 1666464484
transform 1 0 54992 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_487
timestamp 1666464484
transform 1 0 55888 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_489
timestamp 1666464484
transform 1 0 56112 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_492
timestamp 1666464484
transform 1 0 56448 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_508
timestamp 1666464484
transform 1 0 58240 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_5
timestamp 1666464484
transform 1 0 1904 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_21
timestamp 1666464484
transform 1 0 3696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_29
timestamp 1666464484
transform 1 0 4592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_33
timestamp 1666464484
transform 1 0 5040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_37
timestamp 1666464484
transform 1 0 5488 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_53
timestamp 1666464484
transform 1 0 7280 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_63
timestamp 1666464484
transform 1 0 8400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_83
timestamp 1666464484
transform 1 0 10640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_87
timestamp 1666464484
transform 1 0 11088 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_91
timestamp 1666464484
transform 1 0 11536 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_95
timestamp 1666464484
transform 1 0 11984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_105
timestamp 1666464484
transform 1 0 13104 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_109
timestamp 1666464484
transform 1 0 13552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_117
timestamp 1666464484
transform 1 0 14448 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_121
timestamp 1666464484
transform 1 0 14896 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_127
timestamp 1666464484
transform 1 0 15568 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_146
timestamp 1666464484
transform 1 0 17696 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_149
timestamp 1666464484
transform 1 0 18032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_153
timestamp 1666464484
transform 1 0 18480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_157
timestamp 1666464484
transform 1 0 18928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_171
timestamp 1666464484
transform 1 0 20496 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_203
timestamp 1666464484
transform 1 0 24080 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_211
timestamp 1666464484
transform 1 0 24976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_247
timestamp 1666464484
transform 1 0 29008 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_251
timestamp 1666464484
transform 1 0 29456 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_255
timestamp 1666464484
transform 1 0 29904 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_263
timestamp 1666464484
transform 1 0 30800 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_267
timestamp 1666464484
transform 1 0 31248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_271
timestamp 1666464484
transform 1 0 31696 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_275
timestamp 1666464484
transform 1 0 32144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_279
timestamp 1666464484
transform 1 0 32592 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_303
timestamp 1666464484
transform 1 0 35280 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_310
timestamp 1666464484
transform 1 0 36064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_314
timestamp 1666464484
transform 1 0 36512 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_322
timestamp 1666464484
transform 1 0 37408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_326
timestamp 1666464484
transform 1 0 37856 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_328
timestamp 1666464484
transform 1 0 38080 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_331
timestamp 1666464484
transform 1 0 38416 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_335
timestamp 1666464484
transform 1 0 38864 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_351
timestamp 1666464484
transform 1 0 40656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_363
timestamp 1666464484
transform 1 0 42000 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_379
timestamp 1666464484
transform 1 0 43792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_389
timestamp 1666464484
transform 1 0 44912 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_393
timestamp 1666464484
transform 1 0 45360 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_407
timestamp 1666464484
transform 1 0 46928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_411
timestamp 1666464484
transform 1 0 47376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_419
timestamp 1666464484
transform 1 0 48272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_423
timestamp 1666464484
transform 1 0 48720 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1666464484
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_428
timestamp 1666464484
transform 1 0 49280 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_437
timestamp 1666464484
transform 1 0 50288 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_449
timestamp 1666464484
transform 1 0 51632 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_453
timestamp 1666464484
transform 1 0 52080 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_485
timestamp 1666464484
transform 1 0 55664 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_493
timestamp 1666464484
transform 1 0 56560 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_499
timestamp 1666464484
transform 1 0 57232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1666464484
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_9
timestamp 1666464484
transform 1 0 2352 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_17
timestamp 1666464484
transform 1 0 3248 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_33
timestamp 1666464484
transform 1 0 5040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_40
timestamp 1666464484
transform 1 0 5824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_46
timestamp 1666464484
transform 1 0 6496 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_50
timestamp 1666464484
transform 1 0 6944 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_64
timestamp 1666464484
transform 1 0 8512 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_72
timestamp 1666464484
transform 1 0 9408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_76
timestamp 1666464484
transform 1 0 9856 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_80
timestamp 1666464484
transform 1 0 10304 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_84
timestamp 1666464484
transform 1 0 10752 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_88
timestamp 1666464484
transform 1 0 11200 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_91
timestamp 1666464484
transform 1 0 11536 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_108
timestamp 1666464484
transform 1 0 13440 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_121
timestamp 1666464484
transform 1 0 14896 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_127
timestamp 1666464484
transform 1 0 15568 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_135
timestamp 1666464484
transform 1 0 16464 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_141
timestamp 1666464484
transform 1 0 17136 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_145
timestamp 1666464484
transform 1 0 17584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_149
timestamp 1666464484
transform 1 0 18032 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_153
timestamp 1666464484
transform 1 0 18480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_167
timestamp 1666464484
transform 1 0 20048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_171
timestamp 1666464484
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_175
timestamp 1666464484
transform 1 0 20944 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_179
timestamp 1666464484
transform 1 0 21392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_187
timestamp 1666464484
transform 1 0 22288 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_191
timestamp 1666464484
transform 1 0 22736 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 23072 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_200
timestamp 1666464484
transform 1 0 23744 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_202
timestamp 1666464484
transform 1 0 23968 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_205
timestamp 1666464484
transform 1 0 24304 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_219
timestamp 1666464484
transform 1 0 25872 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_223
timestamp 1666464484
transform 1 0 26320 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_227
timestamp 1666464484
transform 1 0 26768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_231
timestamp 1666464484
transform 1 0 27216 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_250
timestamp 1666464484
transform 1 0 29344 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_252
timestamp 1666464484
transform 1 0 29568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_255
timestamp 1666464484
transform 1 0 29904 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_269
timestamp 1666464484
transform 1 0 31472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_273
timestamp 1666464484
transform 1 0 31920 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_278
timestamp 1666464484
transform 1 0 32480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_282
timestamp 1666464484
transform 1 0 32928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_286
timestamp 1666464484
transform 1 0 33376 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_289
timestamp 1666464484
transform 1 0 33712 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_297
timestamp 1666464484
transform 1 0 34608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_301
timestamp 1666464484
transform 1 0 35056 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1666464484
transform 1 0 36848 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_321
timestamp 1666464484
transform 1 0 37296 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_337
timestamp 1666464484
transform 1 0 39088 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_343
timestamp 1666464484
transform 1 0 39760 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_347
timestamp 1666464484
transform 1 0 40208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_361
timestamp 1666464484
transform 1 0 41776 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_369
timestamp 1666464484
transform 1 0 42672 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_373
timestamp 1666464484
transform 1 0 43120 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_377
timestamp 1666464484
transform 1 0 43568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1666464484
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1666464484
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_392
timestamp 1666464484
transform 1 0 45248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_424
timestamp 1666464484
transform 1 0 48832 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_432
timestamp 1666464484
transform 1 0 49728 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_436
timestamp 1666464484
transform 1 0 50176 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_452
timestamp 1666464484
transform 1 0 51968 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1666464484
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_463
timestamp 1666464484
transform 1 0 53200 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_495
timestamp 1666464484
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_503
timestamp 1666464484
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1666464484
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_2
timestamp 1666464484
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_18
timestamp 1666464484
transform 1 0 3360 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_26
timestamp 1666464484
transform 1 0 4256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_30
timestamp 1666464484
transform 1 0 4704 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_32
timestamp 1666464484
transform 1 0 4928 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_35
timestamp 1666464484
transform 1 0 5264 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_51
timestamp 1666464484
transform 1 0 7056 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_59
timestamp 1666464484
transform 1 0 7952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_63
timestamp 1666464484
transform 1 0 8400 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_65
timestamp 1666464484
transform 1 0 8624 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_68
timestamp 1666464484
transform 1 0 8960 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1666464484
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_73
timestamp 1666464484
transform 1 0 9520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_81
timestamp 1666464484
transform 1 0 10416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_87
timestamp 1666464484
transform 1 0 11088 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_91
timestamp 1666464484
transform 1 0 11536 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_97
timestamp 1666464484
transform 1 0 12208 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_111
timestamp 1666464484
transform 1 0 13776 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_115
timestamp 1666464484
transform 1 0 14224 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_119
timestamp 1666464484
transform 1 0 14672 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_123
timestamp 1666464484
transform 1 0 15120 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_127
timestamp 1666464484
transform 1 0 15568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_137
timestamp 1666464484
transform 1 0 16688 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1666464484
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1666464484
transform 1 0 17472 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_149
timestamp 1666464484
transform 1 0 18032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_155
timestamp 1666464484
transform 1 0 18704 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 20272 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_173
timestamp 1666464484
transform 1 0 20720 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_177
timestamp 1666464484
transform 1 0 21168 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_209
timestamp 1666464484
transform 1 0 24752 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1666464484
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1666464484
transform 1 0 25424 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_220
timestamp 1666464484
transform 1 0 25984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_224
timestamp 1666464484
transform 1 0 26432 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_227
timestamp 1666464484
transform 1 0 26768 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_266
timestamp 1666464484
transform 1 0 31136 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_270
timestamp 1666464484
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_278
timestamp 1666464484
transform 1 0 32480 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 32816 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1666464484
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_286
timestamp 1666464484
transform 1 0 33376 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_302
timestamp 1666464484
transform 1 0 35168 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_310
timestamp 1666464484
transform 1 0 36064 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_313
timestamp 1666464484
transform 1 0 36400 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_329
timestamp 1666464484
transform 1 0 38192 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_337
timestamp 1666464484
transform 1 0 39088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_341
timestamp 1666464484
transform 1 0 39536 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_345
timestamp 1666464484
transform 1 0 39984 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1666464484
transform 1 0 40880 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1666464484
transform 1 0 41328 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_360
timestamp 1666464484
transform 1 0 41664 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_424
timestamp 1666464484
transform 1 0 48832 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_428
timestamp 1666464484
transform 1 0 49280 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_441
timestamp 1666464484
transform 1 0 50736 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_445
timestamp 1666464484
transform 1 0 51184 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_477
timestamp 1666464484
transform 1 0 54768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_493
timestamp 1666464484
transform 1 0 56560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_499
timestamp 1666464484
transform 1 0 57232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_507
timestamp 1666464484
transform 1 0 58128 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1666464484
transform 1 0 1568 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_5
timestamp 1666464484
transform 1 0 1904 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_21
timestamp 1666464484
transform 1 0 3696 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_29
timestamp 1666464484
transform 1 0 4592 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_33
timestamp 1666464484
transform 1 0 5040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_37
timestamp 1666464484
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_69
timestamp 1666464484
transform 1 0 9072 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_85
timestamp 1666464484
transform 1 0 10864 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_93
timestamp 1666464484
transform 1 0 11760 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_97
timestamp 1666464484
transform 1 0 12208 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1666464484
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_108
timestamp 1666464484
transform 1 0 13440 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_119
timestamp 1666464484
transform 1 0 14672 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_125
timestamp 1666464484
transform 1 0 15344 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_129
timestamp 1666464484
transform 1 0 15792 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_145
timestamp 1666464484
transform 1 0 17584 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_155
timestamp 1666464484
transform 1 0 18704 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_159
timestamp 1666464484
transform 1 0 19152 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_175
timestamp 1666464484
transform 1 0 20944 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_179
timestamp 1666464484
transform 1 0 21392 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_195
timestamp 1666464484
transform 1 0 23184 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_205
timestamp 1666464484
transform 1 0 24304 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_209
timestamp 1666464484
transform 1 0 24752 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_213
timestamp 1666464484
transform 1 0 25200 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_226
timestamp 1666464484
transform 1 0 26656 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_230
timestamp 1666464484
transform 1 0 27104 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_234
timestamp 1666464484
transform 1 0 27552 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_242
timestamp 1666464484
transform 1 0 28448 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_246
timestamp 1666464484
transform 1 0 28896 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_250
timestamp 1666464484
transform 1 0 29344 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_254
timestamp 1666464484
transform 1 0 29792 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_264
timestamp 1666464484
transform 1 0 30912 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_271
timestamp 1666464484
transform 1 0 31696 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_275
timestamp 1666464484
transform 1 0 32144 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_279
timestamp 1666464484
transform 1 0 32592 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_288
timestamp 1666464484
transform 1 0 33600 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_290
timestamp 1666464484
transform 1 0 33824 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_293
timestamp 1666464484
transform 1 0 34160 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_297
timestamp 1666464484
transform 1 0 34608 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_311
timestamp 1666464484
transform 1 0 36176 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_317
timestamp 1666464484
transform 1 0 36848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_321
timestamp 1666464484
transform 1 0 37296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_329
timestamp 1666464484
transform 1 0 38192 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_333
timestamp 1666464484
transform 1 0 38640 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_335
timestamp 1666464484
transform 1 0 38864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_344
timestamp 1666464484
transform 1 0 39872 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_358
timestamp 1666464484
transform 1 0 41440 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_362
timestamp 1666464484
transform 1 0 41888 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_366
timestamp 1666464484
transform 1 0 42336 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_382
timestamp 1666464484
transform 1 0 44128 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1666464484
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1666464484
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1666464484
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_463
timestamp 1666464484
transform 1 0 53200 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_495
timestamp 1666464484
transform 1 0 56784 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_497
timestamp 1666464484
transform 1 0 57008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_500
timestamp 1666464484
transform 1 0 57344 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_508
timestamp 1666464484
transform 1 0 58240 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1666464484
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_9
timestamp 1666464484
transform 1 0 2352 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_17
timestamp 1666464484
transform 1 0 3248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_25
timestamp 1666464484
transform 1 0 4144 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_29
timestamp 1666464484
transform 1 0 4592 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_61
timestamp 1666464484
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_69
timestamp 1666464484
transform 1 0 9072 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_73
timestamp 1666464484
transform 1 0 9520 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_107
timestamp 1666464484
transform 1 0 13328 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_109
timestamp 1666464484
transform 1 0 13552 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_112
timestamp 1666464484
transform 1 0 13888 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_116
timestamp 1666464484
transform 1 0 14336 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_118
timestamp 1666464484
transform 1 0 14560 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_121
timestamp 1666464484
transform 1 0 14896 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_125
timestamp 1666464484
transform 1 0 15344 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1666464484
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_144
timestamp 1666464484
transform 1 0 17472 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_160
timestamp 1666464484
transform 1 0 19264 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_168
timestamp 1666464484
transform 1 0 20160 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_172
timestamp 1666464484
transform 1 0 20608 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_204
timestamp 1666464484
transform 1 0 24192 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_215
timestamp 1666464484
transform 1 0 25424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_223
timestamp 1666464484
transform 1 0 26320 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_231
timestamp 1666464484
transform 1 0 27216 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_235
timestamp 1666464484
transform 1 0 27664 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_251
timestamp 1666464484
transform 1 0 29456 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_259
timestamp 1666464484
transform 1 0 30352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_263
timestamp 1666464484
transform 1 0 30800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_266
timestamp 1666464484
transform 1 0 31136 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_282
timestamp 1666464484
transform 1 0 32928 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_286
timestamp 1666464484
transform 1 0 33376 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_294
timestamp 1666464484
transform 1 0 34272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_297
timestamp 1666464484
transform 1 0 34608 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_301
timestamp 1666464484
transform 1 0 35056 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_305
timestamp 1666464484
transform 1 0 35504 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_309
timestamp 1666464484
transform 1 0 35952 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_311
timestamp 1666464484
transform 1 0 36176 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_314
timestamp 1666464484
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_330
timestamp 1666464484
transform 1 0 38304 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_333
timestamp 1666464484
transform 1 0 38640 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_353
timestamp 1666464484
transform 1 0 40880 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_357
timestamp 1666464484
transform 1 0 41328 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_360
timestamp 1666464484
transform 1 0 41664 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_364
timestamp 1666464484
transform 1 0 42112 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_380
timestamp 1666464484
transform 1 0 43904 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_384
timestamp 1666464484
transform 1 0 44352 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_388
timestamp 1666464484
transform 1 0 44800 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_402
timestamp 1666464484
transform 1 0 46368 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_406
timestamp 1666464484
transform 1 0 46816 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_422
timestamp 1666464484
transform 1 0 48608 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_428
timestamp 1666464484
transform 1 0 49280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_436
timestamp 1666464484
transform 1 0 50176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_444
timestamp 1666464484
transform 1 0 51072 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_448
timestamp 1666464484
transform 1 0 51520 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_480
timestamp 1666464484
transform 1 0 55104 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1666464484
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1666464484
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1666464484
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1666464484
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1666464484
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1666464484
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1666464484
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1666464484
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_108
timestamp 1666464484
transform 1 0 13440 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_124
timestamp 1666464484
transform 1 0 15232 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_132
timestamp 1666464484
transform 1 0 16128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_168
timestamp 1666464484
transform 1 0 20160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_174
timestamp 1666464484
transform 1 0 20832 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1666464484
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1666464484
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_182
timestamp 1666464484
transform 1 0 21728 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_214
timestamp 1666464484
transform 1 0 25312 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_222
timestamp 1666464484
transform 1 0 26208 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_225
timestamp 1666464484
transform 1 0 26544 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_229
timestamp 1666464484
transform 1 0 26992 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_233
timestamp 1666464484
transform 1 0 27440 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_237
timestamp 1666464484
transform 1 0 27888 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1666464484
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_250
timestamp 1666464484
transform 1 0 29344 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_274
timestamp 1666464484
transform 1 0 32032 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_278
timestamp 1666464484
transform 1 0 32480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_282
timestamp 1666464484
transform 1 0 32928 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_286
timestamp 1666464484
transform 1 0 33376 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_292
timestamp 1666464484
transform 1 0 34048 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_296
timestamp 1666464484
transform 1 0 34496 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_302
timestamp 1666464484
transform 1 0 35168 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_313
timestamp 1666464484
transform 1 0 36400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_317
timestamp 1666464484
transform 1 0 36848 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1666464484
transform 1 0 37296 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_324
timestamp 1666464484
transform 1 0 37632 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_336
timestamp 1666464484
transform 1 0 38976 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_340
timestamp 1666464484
transform 1 0 39424 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_346
timestamp 1666464484
transform 1 0 40096 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_353
timestamp 1666464484
transform 1 0 40880 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_357
timestamp 1666464484
transform 1 0 41328 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_361
timestamp 1666464484
transform 1 0 41776 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_365
timestamp 1666464484
transform 1 0 42224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_369
timestamp 1666464484
transform 1 0 42672 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1666464484
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1666464484
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_392
timestamp 1666464484
transform 1 0 45248 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_400
timestamp 1666464484
transform 1 0 46144 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_404
timestamp 1666464484
transform 1 0 46592 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_407
timestamp 1666464484
transform 1 0 46928 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_417
timestamp 1666464484
transform 1 0 48048 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_427
timestamp 1666464484
transform 1 0 49168 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_431
timestamp 1666464484
transform 1 0 49616 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_447
timestamp 1666464484
transform 1 0 51408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_455
timestamp 1666464484
transform 1 0 52304 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_459
timestamp 1666464484
transform 1 0 52752 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_463
timestamp 1666464484
transform 1 0 53200 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_495
timestamp 1666464484
transform 1 0 56784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_503
timestamp 1666464484
transform 1 0 57680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_507
timestamp 1666464484
transform 1 0 58128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1666464484
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1666464484
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1666464484
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_73
timestamp 1666464484
transform 1 0 9520 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_83
timestamp 1666464484
transform 1 0 10640 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_115
timestamp 1666464484
transform 1 0 14224 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_131
timestamp 1666464484
transform 1 0 16016 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_139
timestamp 1666464484
transform 1 0 16912 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1666464484
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_144
timestamp 1666464484
transform 1 0 17472 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_152
timestamp 1666464484
transform 1 0 18368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_156
timestamp 1666464484
transform 1 0 18816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_192
timestamp 1666464484
transform 1 0 22848 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_196
timestamp 1666464484
transform 1 0 23296 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_200
timestamp 1666464484
transform 1 0 23744 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1666464484
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1666464484
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_215
timestamp 1666464484
transform 1 0 25424 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_221
timestamp 1666464484
transform 1 0 26096 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_225
timestamp 1666464484
transform 1 0 26544 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_229
timestamp 1666464484
transform 1 0 26992 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_242
timestamp 1666464484
transform 1 0 28448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_250
timestamp 1666464484
transform 1 0 29344 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_254
timestamp 1666464484
transform 1 0 29792 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_258
timestamp 1666464484
transform 1 0 30240 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_262
timestamp 1666464484
transform 1 0 30688 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_269
timestamp 1666464484
transform 1 0 31472 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_277
timestamp 1666464484
transform 1 0 32368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 32816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1666464484
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_286
timestamp 1666464484
transform 1 0 33376 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_290
timestamp 1666464484
transform 1 0 33824 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_292
timestamp 1666464484
transform 1 0 34048 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_295
timestamp 1666464484
transform 1 0 34384 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_303
timestamp 1666464484
transform 1 0 35280 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_317
timestamp 1666464484
transform 1 0 36848 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_319
timestamp 1666464484
transform 1 0 37072 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_336
timestamp 1666464484
transform 1 0 38976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_340
timestamp 1666464484
transform 1 0 39424 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_342
timestamp 1666464484
transform 1 0 39648 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_349
timestamp 1666464484
transform 1 0 40432 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_353
timestamp 1666464484
transform 1 0 40880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1666464484
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_360
timestamp 1666464484
transform 1 0 41664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_371
timestamp 1666464484
transform 1 0 42896 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_375
timestamp 1666464484
transform 1 0 43344 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_407
timestamp 1666464484
transform 1 0 46928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_416
timestamp 1666464484
transform 1 0 47936 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_420
timestamp 1666464484
transform 1 0 48384 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_424
timestamp 1666464484
transform 1 0 48832 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1666464484
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1666464484
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1666464484
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_499
timestamp 1666464484
transform 1 0 57232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_507
timestamp 1666464484
transform 1 0 58128 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1666464484
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_5
timestamp 1666464484
transform 1 0 1904 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_21
timestamp 1666464484
transform 1 0 3696 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_29
timestamp 1666464484
transform 1 0 4592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1666464484
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_37
timestamp 1666464484
transform 1 0 5488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_45
timestamp 1666464484
transform 1 0 6384 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_81
timestamp 1666464484
transform 1 0 10416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_87
timestamp 1666464484
transform 1 0 11088 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_91
timestamp 1666464484
transform 1 0 11536 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_99
timestamp 1666464484
transform 1 0 12432 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_103
timestamp 1666464484
transform 1 0 12880 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_108
timestamp 1666464484
transform 1 0 13440 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_174
timestamp 1666464484
transform 1 0 20832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1666464484
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1666464484
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_182
timestamp 1666464484
transform 1 0 21728 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_214
timestamp 1666464484
transform 1 0 25312 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_230
timestamp 1666464484
transform 1 0 27104 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_238
timestamp 1666464484
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_242
timestamp 1666464484
transform 1 0 28448 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_244
timestamp 1666464484
transform 1 0 28672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1666464484
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_250
timestamp 1666464484
transform 1 0 29344 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_257
timestamp 1666464484
transform 1 0 30128 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_273
timestamp 1666464484
transform 1 0 31920 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_281
timestamp 1666464484
transform 1 0 32816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_285
timestamp 1666464484
transform 1 0 33264 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_291
timestamp 1666464484
transform 1 0 33936 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_295
timestamp 1666464484
transform 1 0 34384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_299
timestamp 1666464484
transform 1 0 34832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_303
timestamp 1666464484
transform 1 0 35280 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_307
timestamp 1666464484
transform 1 0 35728 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_311
timestamp 1666464484
transform 1 0 36176 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_315
timestamp 1666464484
transform 1 0 36624 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1666464484
transform 1 0 37296 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_324
timestamp 1666464484
transform 1 0 37632 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_328
timestamp 1666464484
transform 1 0 38080 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_365
timestamp 1666464484
transform 1 0 42224 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_367
timestamp 1666464484
transform 1 0 42448 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_376
timestamp 1666464484
transform 1 0 43456 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_380
timestamp 1666464484
transform 1 0 43904 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_388
timestamp 1666464484
transform 1 0 44800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1666464484
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1666464484
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1666464484
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_463
timestamp 1666464484
transform 1 0 53200 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_495
timestamp 1666464484
transform 1 0 56784 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_497
timestamp 1666464484
transform 1 0 57008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_500
timestamp 1666464484
transform 1 0 57344 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_508
timestamp 1666464484
transform 1 0 58240 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1666464484
transform 1 0 1568 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_9
timestamp 1666464484
transform 1 0 2352 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_41
timestamp 1666464484
transform 1 0 5936 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_57
timestamp 1666464484
transform 1 0 7728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_65
timestamp 1666464484
transform 1 0 8624 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_69
timestamp 1666464484
transform 1 0 9072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_73
timestamp 1666464484
transform 1 0 9520 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_124
timestamp 1666464484
transform 1 0 15232 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_128
timestamp 1666464484
transform 1 0 15680 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_136
timestamp 1666464484
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_140
timestamp 1666464484
transform 1 0 17024 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_144
timestamp 1666464484
transform 1 0 17472 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_160
timestamp 1666464484
transform 1 0 19264 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_162
timestamp 1666464484
transform 1 0 19488 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_165
timestamp 1666464484
transform 1 0 19824 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_201
timestamp 1666464484
transform 1 0 23856 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_205
timestamp 1666464484
transform 1 0 24304 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_209
timestamp 1666464484
transform 1 0 24752 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1666464484
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1666464484
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1666464484
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1666464484
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1666464484
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1666464484
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1666464484
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1666464484
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1666464484
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1666464484
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1666464484
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_499
timestamp 1666464484
transform 1 0 57232 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_507
timestamp 1666464484
transform 1 0 58128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1666464484
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1666464484
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_37
timestamp 1666464484
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_79
timestamp 1666464484
transform 1 0 10192 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_85
timestamp 1666464484
transform 1 0 10864 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_89
timestamp 1666464484
transform 1 0 11312 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_97
timestamp 1666464484
transform 1 0 12208 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_101
timestamp 1666464484
transform 1 0 12656 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1666464484
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1666464484
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_143
timestamp 1666464484
transform 1 0 17360 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_147
timestamp 1666464484
transform 1 0 17808 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_151
timestamp 1666464484
transform 1 0 18256 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_167
timestamp 1666464484
transform 1 0 20048 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_175
timestamp 1666464484
transform 1 0 20944 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1666464484
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1666464484
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1666464484
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_250
timestamp 1666464484
transform 1 0 29344 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_282
timestamp 1666464484
transform 1 0 32928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_286
timestamp 1666464484
transform 1 0 33376 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_299
timestamp 1666464484
transform 1 0 34832 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_307
timestamp 1666464484
transform 1 0 35728 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_313
timestamp 1666464484
transform 1 0 36400 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_317
timestamp 1666464484
transform 1 0 36848 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1666464484
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1666464484
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1666464484
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_392
timestamp 1666464484
transform 1 0 45248 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_397
timestamp 1666464484
transform 1 0 45808 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_401
timestamp 1666464484
transform 1 0 46256 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_433
timestamp 1666464484
transform 1 0 49840 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_449
timestamp 1666464484
transform 1 0 51632 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_457
timestamp 1666464484
transform 1 0 52528 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_463
timestamp 1666464484
transform 1 0 53200 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_495
timestamp 1666464484
transform 1 0 56784 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_503
timestamp 1666464484
transform 1 0 57680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_507
timestamp 1666464484
transform 1 0 58128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_2
timestamp 1666464484
transform 1 0 1568 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_34
timestamp 1666464484
transform 1 0 5152 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1666464484
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_73
timestamp 1666464484
transform 1 0 9520 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_76
timestamp 1666464484
transform 1 0 9856 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_78
timestamp 1666464484
transform 1 0 10080 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_81
timestamp 1666464484
transform 1 0 10416 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_85
timestamp 1666464484
transform 1 0 10864 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_87
timestamp 1666464484
transform 1 0 11088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_90
timestamp 1666464484
transform 1 0 11424 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_94
timestamp 1666464484
transform 1 0 11872 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_98
timestamp 1666464484
transform 1 0 12320 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_102
timestamp 1666464484
transform 1 0 12768 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_138
timestamp 1666464484
transform 1 0 16800 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1666464484
transform 1 0 17472 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_147
timestamp 1666464484
transform 1 0 17808 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_163
timestamp 1666464484
transform 1 0 19600 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_167
timestamp 1666464484
transform 1 0 20048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_203
timestamp 1666464484
transform 1 0 24080 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_207
timestamp 1666464484
transform 1 0 24528 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_211
timestamp 1666464484
transform 1 0 24976 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_215
timestamp 1666464484
transform 1 0 25424 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_247
timestamp 1666464484
transform 1 0 29008 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_255
timestamp 1666464484
transform 1 0 29904 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_259
timestamp 1666464484
transform 1 0 30352 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_262
timestamp 1666464484
transform 1 0 30688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_266
timestamp 1666464484
transform 1 0 31136 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_272
timestamp 1666464484
transform 1 0 31808 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_276
timestamp 1666464484
transform 1 0 32256 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_280
timestamp 1666464484
transform 1 0 32704 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_286
timestamp 1666464484
transform 1 0 33376 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_288
timestamp 1666464484
transform 1 0 33600 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_293
timestamp 1666464484
transform 1 0 34160 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_303
timestamp 1666464484
transform 1 0 35280 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_307
timestamp 1666464484
transform 1 0 35728 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_311
timestamp 1666464484
transform 1 0 36176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_325
timestamp 1666464484
transform 1 0 37744 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_341
timestamp 1666464484
transform 1 0 39536 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_349
timestamp 1666464484
transform 1 0 40432 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_353
timestamp 1666464484
transform 1 0 40880 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1666464484
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_421
timestamp 1666464484
transform 1 0 48496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1666464484
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1666464484
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1666464484
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1666464484
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_499
timestamp 1666464484
transform 1 0 57232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_507
timestamp 1666464484
transform 1 0 58128 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1666464484
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_5
timestamp 1666464484
transform 1 0 1904 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_21
timestamp 1666464484
transform 1 0 3696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_29
timestamp 1666464484
transform 1 0 4592 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1666464484
transform 1 0 5040 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_37
timestamp 1666464484
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_53
timestamp 1666464484
transform 1 0 7280 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_88
timestamp 1666464484
transform 1 0 11200 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_94
timestamp 1666464484
transform 1 0 11872 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_98
timestamp 1666464484
transform 1 0 12320 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_108
timestamp 1666464484
transform 1 0 13440 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_118
timestamp 1666464484
transform 1 0 14560 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_154
timestamp 1666464484
transform 1 0 18592 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_158
timestamp 1666464484
transform 1 0 19040 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_162
timestamp 1666464484
transform 1 0 19488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_170
timestamp 1666464484
transform 1 0 20384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_174
timestamp 1666464484
transform 1 0 20832 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1666464484
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1666464484
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_243
timestamp 1666464484
transform 1 0 28560 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1666464484
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_250
timestamp 1666464484
transform 1 0 29344 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_254
timestamp 1666464484
transform 1 0 29792 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_260
timestamp 1666464484
transform 1 0 30464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_268
timestamp 1666464484
transform 1 0 31360 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_270
timestamp 1666464484
transform 1 0 31584 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_275
timestamp 1666464484
transform 1 0 32144 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_281
timestamp 1666464484
transform 1 0 32816 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_285
timestamp 1666464484
transform 1 0 33264 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_289
timestamp 1666464484
transform 1 0 33712 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_305
timestamp 1666464484
transform 1 0 35504 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_313
timestamp 1666464484
transform 1 0 36400 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_317
timestamp 1666464484
transform 1 0 36848 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_321
timestamp 1666464484
transform 1 0 37296 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_337
timestamp 1666464484
transform 1 0 39088 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_345
timestamp 1666464484
transform 1 0 39984 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_349
timestamp 1666464484
transform 1 0 40432 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_381
timestamp 1666464484
transform 1 0 44016 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1666464484
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1666464484
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_456
timestamp 1666464484
transform 1 0 52416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1666464484
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_463
timestamp 1666464484
transform 1 0 53200 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_495
timestamp 1666464484
transform 1 0 56784 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_497
timestamp 1666464484
transform 1 0 57008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_500
timestamp 1666464484
transform 1 0 57344 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_508
timestamp 1666464484
transform 1 0 58240 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1666464484
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_9
timestamp 1666464484
transform 1 0 2352 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_25
timestamp 1666464484
transform 1 0 4144 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_33
timestamp 1666464484
transform 1 0 5040 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_35
timestamp 1666464484
transform 1 0 5264 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1666464484
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1666464484
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_76
timestamp 1666464484
transform 1 0 9856 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_80
timestamp 1666464484
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_86
timestamp 1666464484
transform 1 0 10976 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_90
timestamp 1666464484
transform 1 0 11424 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_122
timestamp 1666464484
transform 1 0 15008 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_138
timestamp 1666464484
transform 1 0 16800 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_144
timestamp 1666464484
transform 1 0 17472 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_160
timestamp 1666464484
transform 1 0 19264 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 19936 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_202
timestamp 1666464484
transform 1 0 23968 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_206
timestamp 1666464484
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_210
timestamp 1666464484
transform 1 0 24864 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1666464484
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_215
timestamp 1666464484
transform 1 0 25424 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_231
timestamp 1666464484
transform 1 0 27216 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_235
timestamp 1666464484
transform 1 0 27664 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_239
timestamp 1666464484
transform 1 0 28112 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_245
timestamp 1666464484
transform 1 0 28784 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_247
timestamp 1666464484
transform 1 0 29008 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_260
timestamp 1666464484
transform 1 0 30464 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_264
timestamp 1666464484
transform 1 0 30912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_266
timestamp 1666464484
transform 1 0 31136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_271
timestamp 1666464484
transform 1 0 31696 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_277
timestamp 1666464484
transform 1 0 32368 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 32816 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1666464484
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_286
timestamp 1666464484
transform 1 0 33376 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_302
timestamp 1666464484
transform 1 0 35168 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_310
timestamp 1666464484
transform 1 0 36064 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_314
timestamp 1666464484
transform 1 0 36512 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_316
timestamp 1666464484
transform 1 0 36736 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_323
timestamp 1666464484
transform 1 0 37520 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_327
timestamp 1666464484
transform 1 0 37968 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_331
timestamp 1666464484
transform 1 0 38416 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_339
timestamp 1666464484
transform 1 0 39312 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_347
timestamp 1666464484
transform 1 0 40208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_349
timestamp 1666464484
transform 1 0 40432 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1666464484
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_357
timestamp 1666464484
transform 1 0 41328 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_360
timestamp 1666464484
transform 1 0 41664 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_424
timestamp 1666464484
transform 1 0 48832 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1666464484
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1666464484
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1666464484
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_499
timestamp 1666464484
transform 1 0 57232 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_507
timestamp 1666464484
transform 1 0 58128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1666464484
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1666464484
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_37
timestamp 1666464484
transform 1 0 5488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_45
timestamp 1666464484
transform 1 0 6384 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_49
timestamp 1666464484
transform 1 0 6832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_84
timestamp 1666464484
transform 1 0 10752 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_90
timestamp 1666464484
transform 1 0 11424 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_94
timestamp 1666464484
transform 1 0 11872 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_102
timestamp 1666464484
transform 1 0 12768 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_108
timestamp 1666464484
transform 1 0 13440 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_124
timestamp 1666464484
transform 1 0 15232 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_166
timestamp 1666464484
transform 1 0 19936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_172
timestamp 1666464484
transform 1 0 20608 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1666464484
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1666464484
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_243
timestamp 1666464484
transform 1 0 28560 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_246
timestamp 1666464484
transform 1 0 28896 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_250
timestamp 1666464484
transform 1 0 29344 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_258
timestamp 1666464484
transform 1 0 30240 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_264
timestamp 1666464484
transform 1 0 30912 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_268
timestamp 1666464484
transform 1 0 31360 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_270
timestamp 1666464484
transform 1 0 31584 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_273
timestamp 1666464484
transform 1 0 31920 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_279
timestamp 1666464484
transform 1 0 32592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_287
timestamp 1666464484
transform 1 0 33488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_289
timestamp 1666464484
transform 1 0 33712 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_294
timestamp 1666464484
transform 1 0 34272 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_298
timestamp 1666464484
transform 1 0 34720 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_302
timestamp 1666464484
transform 1 0 35168 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_305
timestamp 1666464484
transform 1 0 35504 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_313
timestamp 1666464484
transform 1 0 36400 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_317
timestamp 1666464484
transform 1 0 36848 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1666464484
transform 1 0 37296 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_334
timestamp 1666464484
transform 1 0 38752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_338
timestamp 1666464484
transform 1 0 39200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_346
timestamp 1666464484
transform 1 0 40096 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_350
timestamp 1666464484
transform 1 0 40544 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_382
timestamp 1666464484
transform 1 0 44128 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1666464484
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1666464484
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1666464484
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_463
timestamp 1666464484
transform 1 0 53200 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_495
timestamp 1666464484
transform 1 0 56784 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_503
timestamp 1666464484
transform 1 0 57680 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_507
timestamp 1666464484
transform 1 0 58128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_2
timestamp 1666464484
transform 1 0 1568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_10
timestamp 1666464484
transform 1 0 2464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_14
timestamp 1666464484
transform 1 0 2912 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_18
timestamp 1666464484
transform 1 0 3360 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_26
timestamp 1666464484
transform 1 0 4256 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_30
timestamp 1666464484
transform 1 0 4704 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_62
timestamp 1666464484
transform 1 0 8288 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1666464484
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_73
timestamp 1666464484
transform 1 0 9520 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_76
timestamp 1666464484
transform 1 0 9856 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_92
timestamp 1666464484
transform 1 0 11648 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_96
timestamp 1666464484
transform 1 0 12096 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_100
timestamp 1666464484
transform 1 0 12544 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_132
timestamp 1666464484
transform 1 0 16128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_140
timestamp 1666464484
transform 1 0 17024 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_144
timestamp 1666464484
transform 1 0 17472 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_160
timestamp 1666464484
transform 1 0 19264 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_164
timestamp 1666464484
transform 1 0 19712 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_168
timestamp 1666464484
transform 1 0 20160 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_204
timestamp 1666464484
transform 1 0 24192 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1666464484
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1666464484
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_215
timestamp 1666464484
transform 1 0 25424 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_231
timestamp 1666464484
transform 1 0 27216 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_233
timestamp 1666464484
transform 1 0 27440 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_238
timestamp 1666464484
transform 1 0 28000 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_242
timestamp 1666464484
transform 1 0 28448 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_246
timestamp 1666464484
transform 1 0 28896 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_248
timestamp 1666464484
transform 1 0 29120 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_253
timestamp 1666464484
transform 1 0 29680 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_257
timestamp 1666464484
transform 1 0 30128 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_273
timestamp 1666464484
transform 1 0 31920 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1666464484
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_286
timestamp 1666464484
transform 1 0 33376 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_291
timestamp 1666464484
transform 1 0 33936 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_297
timestamp 1666464484
transform 1 0 34608 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_301
timestamp 1666464484
transform 1 0 35056 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_317
timestamp 1666464484
transform 1 0 36848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_320
timestamp 1666464484
transform 1 0 37184 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_324
timestamp 1666464484
transform 1 0 37632 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_340
timestamp 1666464484
transform 1 0 39424 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_348
timestamp 1666464484
transform 1 0 40320 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_352
timestamp 1666464484
transform 1 0 40768 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1666464484
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_357
timestamp 1666464484
transform 1 0 41328 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_363
timestamp 1666464484
transform 1 0 42000 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_367
timestamp 1666464484
transform 1 0 42448 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_381
timestamp 1666464484
transform 1 0 44016 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_397
timestamp 1666464484
transform 1 0 45808 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_405
timestamp 1666464484
transform 1 0 46704 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_409
timestamp 1666464484
transform 1 0 47152 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_411
timestamp 1666464484
transform 1 0 47376 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_420
timestamp 1666464484
transform 1 0 48384 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_424
timestamp 1666464484
transform 1 0 48832 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1666464484
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1666464484
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1666464484
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_499
timestamp 1666464484
transform 1 0 57232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_507
timestamp 1666464484
transform 1 0 58128 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_2
timestamp 1666464484
transform 1 0 1568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_10
timestamp 1666464484
transform 1 0 2464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_14
timestamp 1666464484
transform 1 0 2912 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_16
timestamp 1666464484
transform 1 0 3136 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_19
timestamp 1666464484
transform 1 0 3472 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_37
timestamp 1666464484
transform 1 0 5488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_53
timestamp 1666464484
transform 1 0 7280 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_61
timestamp 1666464484
transform 1 0 8176 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_96
timestamp 1666464484
transform 1 0 12096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_102
timestamp 1666464484
transform 1 0 12768 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1666464484
transform 1 0 13440 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_159
timestamp 1666464484
transform 1 0 19152 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_163
timestamp 1666464484
transform 1 0 19600 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_171
timestamp 1666464484
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_175
timestamp 1666464484
transform 1 0 20944 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_179
timestamp 1666464484
transform 1 0 21392 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_211
timestamp 1666464484
transform 1 0 24976 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_219
timestamp 1666464484
transform 1 0 25872 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_223
timestamp 1666464484
transform 1 0 26320 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_225
timestamp 1666464484
transform 1 0 26544 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_228
timestamp 1666464484
transform 1 0 26880 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_234
timestamp 1666464484
transform 1 0 27552 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_240
timestamp 1666464484
transform 1 0 28224 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_246
timestamp 1666464484
transform 1 0 28896 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_250
timestamp 1666464484
transform 1 0 29344 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_253
timestamp 1666464484
transform 1 0 29680 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_317
timestamp 1666464484
transform 1 0 36848 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1666464484
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1666464484
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1666464484
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_392
timestamp 1666464484
transform 1 0 45248 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_400
timestamp 1666464484
transform 1 0 46144 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_404
timestamp 1666464484
transform 1 0 46592 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_408
timestamp 1666464484
transform 1 0 47040 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_412
timestamp 1666464484
transform 1 0 47488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_424
timestamp 1666464484
transform 1 0 48832 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_428
timestamp 1666464484
transform 1 0 49280 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1666464484
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_463
timestamp 1666464484
transform 1 0 53200 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_495
timestamp 1666464484
transform 1 0 56784 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_503
timestamp 1666464484
transform 1 0 57680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_507
timestamp 1666464484
transform 1 0 58128 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_2
timestamp 1666464484
transform 1 0 1568 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_17
timestamp 1666464484
transform 1 0 3248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_19
timestamp 1666464484
transform 1 0 3472 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_26
timestamp 1666464484
transform 1 0 4256 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_30
timestamp 1666464484
transform 1 0 4704 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_62
timestamp 1666464484
transform 1 0 8288 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1666464484
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_73
timestamp 1666464484
transform 1 0 9520 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_83
timestamp 1666464484
transform 1 0 10640 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_91
timestamp 1666464484
transform 1 0 11536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_95
timestamp 1666464484
transform 1 0 11984 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_98
timestamp 1666464484
transform 1 0 12320 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_130
timestamp 1666464484
transform 1 0 15904 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_138
timestamp 1666464484
transform 1 0 16800 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1666464484
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1666464484
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1666464484
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_215
timestamp 1666464484
transform 1 0 25424 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_231
timestamp 1666464484
transform 1 0 27216 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_237
timestamp 1666464484
transform 1 0 27888 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_241
timestamp 1666464484
transform 1 0 28336 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_246
timestamp 1666464484
transform 1 0 28896 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_250
timestamp 1666464484
transform 1 0 29344 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_282
timestamp 1666464484
transform 1 0 32928 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_286
timestamp 1666464484
transform 1 0 33376 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_318
timestamp 1666464484
transform 1 0 36960 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_322
timestamp 1666464484
transform 1 0 37408 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_324
timestamp 1666464484
transform 1 0 37632 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_329
timestamp 1666464484
transform 1 0 38192 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_333
timestamp 1666464484
transform 1 0 38640 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_349
timestamp 1666464484
transform 1 0 40432 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_353
timestamp 1666464484
transform 1 0 40880 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_357
timestamp 1666464484
transform 1 0 41328 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_389
timestamp 1666464484
transform 1 0 44912 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_397
timestamp 1666464484
transform 1 0 45808 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_401
timestamp 1666464484
transform 1 0 46256 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_403
timestamp 1666464484
transform 1 0 46480 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_406
timestamp 1666464484
transform 1 0 46816 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_410
timestamp 1666464484
transform 1 0 47264 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_424
timestamp 1666464484
transform 1 0 48832 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1666464484
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1666464484
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1666464484
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_499
timestamp 1666464484
transform 1 0 57232 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_507
timestamp 1666464484
transform 1 0 58128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1666464484
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1666464484
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_37
timestamp 1666464484
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_45
timestamp 1666464484
transform 1 0 6384 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_81
timestamp 1666464484
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_87
timestamp 1666464484
transform 1 0 11088 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_91
timestamp 1666464484
transform 1 0 11536 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_99
timestamp 1666464484
transform 1 0 12432 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_103
timestamp 1666464484
transform 1 0 12880 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1666464484
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_108
timestamp 1666464484
transform 1 0 13440 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_174
timestamp 1666464484
transform 1 0 20832 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1666464484
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_179
timestamp 1666464484
transform 1 0 21392 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_182
timestamp 1666464484
transform 1 0 21728 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_214
timestamp 1666464484
transform 1 0 25312 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_230
timestamp 1666464484
transform 1 0 27104 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_234
timestamp 1666464484
transform 1 0 27552 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_236
timestamp 1666464484
transform 1 0 27776 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_239
timestamp 1666464484
transform 1 0 28112 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1666464484
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_250
timestamp 1666464484
transform 1 0 29344 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_266
timestamp 1666464484
transform 1 0 31136 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_270
timestamp 1666464484
transform 1 0 31584 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_275
timestamp 1666464484
transform 1 0 32144 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_279
timestamp 1666464484
transform 1 0 32592 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_295
timestamp 1666464484
transform 1 0 34384 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_303
timestamp 1666464484
transform 1 0 35280 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_315
timestamp 1666464484
transform 1 0 36624 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1666464484
transform 1 0 37296 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_324
timestamp 1666464484
transform 1 0 37632 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_388
timestamp 1666464484
transform 1 0 44800 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_392
timestamp 1666464484
transform 1 0 45248 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_408
timestamp 1666464484
transform 1 0 47040 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_414
timestamp 1666464484
transform 1 0 47712 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_446
timestamp 1666464484
transform 1 0 51296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_454
timestamp 1666464484
transform 1 0 52192 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_458
timestamp 1666464484
transform 1 0 52640 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1666464484
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_463
timestamp 1666464484
transform 1 0 53200 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_495
timestamp 1666464484
transform 1 0 56784 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_503
timestamp 1666464484
transform 1 0 57680 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_507
timestamp 1666464484
transform 1 0 58128 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_2
timestamp 1666464484
transform 1 0 1568 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_5
timestamp 1666464484
transform 1 0 1904 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_69
timestamp 1666464484
transform 1 0 9072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_73
timestamp 1666464484
transform 1 0 9520 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_124
timestamp 1666464484
transform 1 0 15232 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_128
timestamp 1666464484
transform 1 0 15680 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_136
timestamp 1666464484
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_140
timestamp 1666464484
transform 1 0 17024 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_144
timestamp 1666464484
transform 1 0 17472 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_152
timestamp 1666464484
transform 1 0 18368 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_155
timestamp 1666464484
transform 1 0 18704 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_191
timestamp 1666464484
transform 1 0 22736 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_195
timestamp 1666464484
transform 1 0 23184 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_211
timestamp 1666464484
transform 1 0 24976 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_215
timestamp 1666464484
transform 1 0 25424 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_247
timestamp 1666464484
transform 1 0 29008 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_263
timestamp 1666464484
transform 1 0 30800 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_271
timestamp 1666464484
transform 1 0 31696 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_277
timestamp 1666464484
transform 1 0 32368 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_281
timestamp 1666464484
transform 1 0 32816 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1666464484
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_286
timestamp 1666464484
transform 1 0 33376 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_302
timestamp 1666464484
transform 1 0 35168 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_306
timestamp 1666464484
transform 1 0 35616 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_315
timestamp 1666464484
transform 1 0 36624 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_319
timestamp 1666464484
transform 1 0 37072 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_351
timestamp 1666464484
transform 1 0 40656 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_357
timestamp 1666464484
transform 1 0 41328 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_373
timestamp 1666464484
transform 1 0 43120 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_379
timestamp 1666464484
transform 1 0 43792 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_387
timestamp 1666464484
transform 1 0 44688 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_391
timestamp 1666464484
transform 1 0 45136 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_423
timestamp 1666464484
transform 1 0 48720 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1666464484
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1666464484
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1666464484
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1666464484
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_499
timestamp 1666464484
transform 1 0 57232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_507
timestamp 1666464484
transform 1 0 58128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_2
timestamp 1666464484
transform 1 0 1568 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_9
timestamp 1666464484
transform 1 0 2352 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_25
timestamp 1666464484
transform 1 0 4144 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_33
timestamp 1666464484
transform 1 0 5040 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_37
timestamp 1666464484
transform 1 0 5488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_53
timestamp 1666464484
transform 1 0 7280 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_57
timestamp 1666464484
transform 1 0 7728 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_93
timestamp 1666464484
transform 1 0 11760 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_99
timestamp 1666464484
transform 1 0 12432 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_103
timestamp 1666464484
transform 1 0 12880 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1666464484
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_108
timestamp 1666464484
transform 1 0 13440 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_116
timestamp 1666464484
transform 1 0 14336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_120
timestamp 1666464484
transform 1 0 14784 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_155
timestamp 1666464484
transform 1 0 18704 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_161
timestamp 1666464484
transform 1 0 19376 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_165
timestamp 1666464484
transform 1 0 19824 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_173
timestamp 1666464484
transform 1 0 20720 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1666464484
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1666464484
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1666464484
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_250
timestamp 1666464484
transform 1 0 29344 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_266
timestamp 1666464484
transform 1 0 31136 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_274
timestamp 1666464484
transform 1 0 32032 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_276
timestamp 1666464484
transform 1 0 32256 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_279
timestamp 1666464484
transform 1 0 32592 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_295
timestamp 1666464484
transform 1 0 34384 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_303
timestamp 1666464484
transform 1 0 35280 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_312
timestamp 1666464484
transform 1 0 36288 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_316
timestamp 1666464484
transform 1 0 36736 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1666464484
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_321
timestamp 1666464484
transform 1 0 37296 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_337
timestamp 1666464484
transform 1 0 39088 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_339
timestamp 1666464484
transform 1 0 39312 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_342
timestamp 1666464484
transform 1 0 39648 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_344
timestamp 1666464484
transform 1 0 39872 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_351
timestamp 1666464484
transform 1 0 40656 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_355
timestamp 1666464484
transform 1 0 41104 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_387
timestamp 1666464484
transform 1 0 44688 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1666464484
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1666464484
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1666464484
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1666464484
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_463
timestamp 1666464484
transform 1 0 53200 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_495
timestamp 1666464484
transform 1 0 56784 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_497
timestamp 1666464484
transform 1 0 57008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_500
timestamp 1666464484
transform 1 0 57344 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_508
timestamp 1666464484
transform 1 0 58240 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_2
timestamp 1666464484
transform 1 0 1568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_18
timestamp 1666464484
transform 1 0 3360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_26
timestamp 1666464484
transform 1 0 4256 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_32
timestamp 1666464484
transform 1 0 4928 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_36
timestamp 1666464484
transform 1 0 5376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_68
timestamp 1666464484
transform 1 0 8960 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1666464484
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_73
timestamp 1666464484
transform 1 0 9520 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_81
timestamp 1666464484
transform 1 0 10416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_85
timestamp 1666464484
transform 1 0 10864 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_88
timestamp 1666464484
transform 1 0 11200 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_92
timestamp 1666464484
transform 1 0 11648 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_95
timestamp 1666464484
transform 1 0 11984 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_127
timestamp 1666464484
transform 1 0 15568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_135
timestamp 1666464484
transform 1 0 16464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_139
timestamp 1666464484
transform 1 0 16912 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1666464484
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_144
timestamp 1666464484
transform 1 0 17472 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_148
timestamp 1666464484
transform 1 0 17920 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_150
timestamp 1666464484
transform 1 0 18144 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_153
timestamp 1666464484
transform 1 0 18480 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_157
timestamp 1666464484
transform 1 0 18928 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_161
timestamp 1666464484
transform 1 0 19376 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_196
timestamp 1666464484
transform 1 0 23296 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_200
timestamp 1666464484
transform 1 0 23744 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1666464484
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1666464484
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1666464484
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1666464484
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1666464484
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_286
timestamp 1666464484
transform 1 0 33376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_318
timestamp 1666464484
transform 1 0 36960 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_326
timestamp 1666464484
transform 1 0 37856 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_330
timestamp 1666464484
transform 1 0 38304 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_334
timestamp 1666464484
transform 1 0 38752 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_338
timestamp 1666464484
transform 1 0 39200 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1666464484
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_357
timestamp 1666464484
transform 1 0 41328 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_360
timestamp 1666464484
transform 1 0 41664 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_362
timestamp 1666464484
transform 1 0 41888 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_365
timestamp 1666464484
transform 1 0 42224 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_369
timestamp 1666464484
transform 1 0 42672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_383
timestamp 1666464484
transform 1 0 44240 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_415
timestamp 1666464484
transform 1 0 47824 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_423
timestamp 1666464484
transform 1 0 48720 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1666464484
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_428
timestamp 1666464484
transform 1 0 49280 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_460
timestamp 1666464484
transform 1 0 52864 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_464
timestamp 1666464484
transform 1 0 53312 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1666464484
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_499
timestamp 1666464484
transform 1 0 57232 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1666464484
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1666464484
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1666464484
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_37
timestamp 1666464484
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_45
timestamp 1666464484
transform 1 0 6384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_49
timestamp 1666464484
transform 1 0 6832 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_51
timestamp 1666464484
transform 1 0 7056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_86
timestamp 1666464484
transform 1 0 10976 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_92
timestamp 1666464484
transform 1 0 11648 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_96
timestamp 1666464484
transform 1 0 12096 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_104
timestamp 1666464484
transform 1 0 12992 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_108
timestamp 1666464484
transform 1 0 13440 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_124
timestamp 1666464484
transform 1 0 15232 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_132
timestamp 1666464484
transform 1 0 16128 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_167
timestamp 1666464484
transform 1 0 20048 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_173
timestamp 1666464484
transform 1 0 20720 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_179
timestamp 1666464484
transform 1 0 21392 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_182
timestamp 1666464484
transform 1 0 21728 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_186
timestamp 1666464484
transform 1 0 22176 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_218
timestamp 1666464484
transform 1 0 25760 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_236
timestamp 1666464484
transform 1 0 27776 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_244
timestamp 1666464484
transform 1 0 28672 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_250
timestamp 1666464484
transform 1 0 29344 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_253
timestamp 1666464484
transform 1 0 29680 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_255
timestamp 1666464484
transform 1 0 29904 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_258
timestamp 1666464484
transform 1 0 30240 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_264
timestamp 1666464484
transform 1 0 30912 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_266
timestamp 1666464484
transform 1 0 31136 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_271
timestamp 1666464484
transform 1 0 31696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_275
timestamp 1666464484
transform 1 0 32144 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_307
timestamp 1666464484
transform 1 0 35728 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_315
timestamp 1666464484
transform 1 0 36624 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1666464484
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1666464484
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1666464484
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_392
timestamp 1666464484
transform 1 0 45248 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_424
timestamp 1666464484
transform 1 0 48832 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_440
timestamp 1666464484
transform 1 0 50624 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_444
timestamp 1666464484
transform 1 0 51072 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_452
timestamp 1666464484
transform 1 0 51968 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_456
timestamp 1666464484
transform 1 0 52416 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1666464484
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_463
timestamp 1666464484
transform 1 0 53200 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_476
timestamp 1666464484
transform 1 0 54656 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_508
timestamp 1666464484
transform 1 0 58240 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1666464484
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_5
timestamp 1666464484
transform 1 0 1904 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_13
timestamp 1666464484
transform 1 0 2800 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_17
timestamp 1666464484
transform 1 0 3248 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_19
timestamp 1666464484
transform 1 0 3472 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_26
timestamp 1666464484
transform 1 0 4256 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_30
timestamp 1666464484
transform 1 0 4704 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_34
timestamp 1666464484
transform 1 0 5152 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1666464484
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_73
timestamp 1666464484
transform 1 0 9520 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_76
timestamp 1666464484
transform 1 0 9856 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_80
timestamp 1666464484
transform 1 0 10304 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_84
timestamp 1666464484
transform 1 0 10752 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_92
timestamp 1666464484
transform 1 0 11648 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_96
timestamp 1666464484
transform 1 0 12096 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_98
timestamp 1666464484
transform 1 0 12320 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_101
timestamp 1666464484
transform 1 0 12656 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_105
timestamp 1666464484
transform 1 0 13104 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1666464484
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_144
timestamp 1666464484
transform 1 0 17472 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_147
timestamp 1666464484
transform 1 0 17808 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_151
timestamp 1666464484
transform 1 0 18256 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_155
timestamp 1666464484
transform 1 0 18704 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_163
timestamp 1666464484
transform 1 0 19600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_165
timestamp 1666464484
transform 1 0 19824 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_168
timestamp 1666464484
transform 1 0 20160 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_204
timestamp 1666464484
transform 1 0 24192 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1666464484
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1666464484
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_215
timestamp 1666464484
transform 1 0 25424 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_223
timestamp 1666464484
transform 1 0 26320 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_227
timestamp 1666464484
transform 1 0 26768 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_229
timestamp 1666464484
transform 1 0 26992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_234
timestamp 1666464484
transform 1 0 27552 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_242
timestamp 1666464484
transform 1 0 28448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_250
timestamp 1666464484
transform 1 0 29344 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_256
timestamp 1666464484
transform 1 0 30016 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_262
timestamp 1666464484
transform 1 0 30688 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_268
timestamp 1666464484
transform 1 0 31360 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_272
timestamp 1666464484
transform 1 0 31808 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_280
timestamp 1666464484
transform 1 0 32704 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_286
timestamp 1666464484
transform 1 0 33376 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_318
timestamp 1666464484
transform 1 0 36960 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_334
timestamp 1666464484
transform 1 0 38752 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_338
timestamp 1666464484
transform 1 0 39200 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_342
timestamp 1666464484
transform 1 0 39648 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_350
timestamp 1666464484
transform 1 0 40544 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1666464484
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_357
timestamp 1666464484
transform 1 0 41328 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_360
timestamp 1666464484
transform 1 0 41664 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_368
timestamp 1666464484
transform 1 0 42560 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_371
timestamp 1666464484
transform 1 0 42896 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_379
timestamp 1666464484
transform 1 0 43792 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_383
timestamp 1666464484
transform 1 0 44240 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_415
timestamp 1666464484
transform 1 0 47824 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_423
timestamp 1666464484
transform 1 0 48720 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1666464484
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1666464484
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1666464484
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1666464484
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1666464484
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_507
timestamp 1666464484
transform 1 0 58128 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1666464484
transform 1 0 1568 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_9
timestamp 1666464484
transform 1 0 2352 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_17
timestamp 1666464484
transform 1 0 3248 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_19
timestamp 1666464484
transform 1 0 3472 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_26
timestamp 1666464484
transform 1 0 4256 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_30
timestamp 1666464484
transform 1 0 4704 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1666464484
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_37
timestamp 1666464484
transform 1 0 5488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_53
timestamp 1666464484
transform 1 0 7280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_61
timestamp 1666464484
transform 1 0 8176 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_97
timestamp 1666464484
transform 1 0 12208 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_103
timestamp 1666464484
transform 1 0 12880 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1666464484
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_108
timestamp 1666464484
transform 1 0 13440 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_110
timestamp 1666464484
transform 1 0 13664 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_113
timestamp 1666464484
transform 1 0 14000 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_149
timestamp 1666464484
transform 1 0 18032 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_153
timestamp 1666464484
transform 1 0 18480 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_157
timestamp 1666464484
transform 1 0 18928 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_173
timestamp 1666464484
transform 1 0 20720 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_179
timestamp 1666464484
transform 1 0 21392 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_211
timestamp 1666464484
transform 1 0 24976 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_227
timestamp 1666464484
transform 1 0 26768 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_235
timestamp 1666464484
transform 1 0 27664 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_241
timestamp 1666464484
transform 1 0 28336 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1666464484
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_250
timestamp 1666464484
transform 1 0 29344 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_253
timestamp 1666464484
transform 1 0 29680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_261
timestamp 1666464484
transform 1 0 30576 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_267
timestamp 1666464484
transform 1 0 31248 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_271
timestamp 1666464484
transform 1 0 31696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_275
timestamp 1666464484
transform 1 0 32144 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_281
timestamp 1666464484
transform 1 0 32816 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_285
timestamp 1666464484
transform 1 0 33264 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_317
timestamp 1666464484
transform 1 0 36848 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_321
timestamp 1666464484
transform 1 0 37296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_329
timestamp 1666464484
transform 1 0 38192 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_332
timestamp 1666464484
transform 1 0 38528 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_340
timestamp 1666464484
transform 1 0 39424 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_348
timestamp 1666464484
transform 1 0 40320 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_352
timestamp 1666464484
transform 1 0 40768 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_368
timestamp 1666464484
transform 1 0 42560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_372
timestamp 1666464484
transform 1 0 43008 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_388
timestamp 1666464484
transform 1 0 44800 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_392
timestamp 1666464484
transform 1 0 45248 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_397
timestamp 1666464484
transform 1 0 45808 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_401
timestamp 1666464484
transform 1 0 46256 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_433
timestamp 1666464484
transform 1 0 49840 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_449
timestamp 1666464484
transform 1 0 51632 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_457
timestamp 1666464484
transform 1 0 52528 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1666464484
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1666464484
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_503
timestamp 1666464484
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_507
timestamp 1666464484
transform 1 0 58128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_2
timestamp 1666464484
transform 1 0 1568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_5
timestamp 1666464484
transform 1 0 1904 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_69
timestamp 1666464484
transform 1 0 9072 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_73
timestamp 1666464484
transform 1 0 9520 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_89
timestamp 1666464484
transform 1 0 11312 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_92
timestamp 1666464484
transform 1 0 11648 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_96
timestamp 1666464484
transform 1 0 12096 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_99
timestamp 1666464484
transform 1 0 12432 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_131
timestamp 1666464484
transform 1 0 16016 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_139
timestamp 1666464484
transform 1 0 16912 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1666464484
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_144
timestamp 1666464484
transform 1 0 17472 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_160
timestamp 1666464484
transform 1 0 19264 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_162
timestamp 1666464484
transform 1 0 19488 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_165
timestamp 1666464484
transform 1 0 19824 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_201
timestamp 1666464484
transform 1 0 23856 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_205
timestamp 1666464484
transform 1 0 24304 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_215
timestamp 1666464484
transform 1 0 25424 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_231
timestamp 1666464484
transform 1 0 27216 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_237
timestamp 1666464484
transform 1 0 27888 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_245
timestamp 1666464484
transform 1 0 28784 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_249
timestamp 1666464484
transform 1 0 29232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_257
timestamp 1666464484
transform 1 0 30128 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_263
timestamp 1666464484
transform 1 0 30800 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1666464484
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1666464484
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1666464484
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1666464484
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1666464484
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1666464484
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1666464484
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1666464484
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1666464484
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1666464484
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1666464484
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_499
timestamp 1666464484
transform 1 0 57232 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 57680 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_508
timestamp 1666464484
transform 1 0 58240 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1666464484
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_9
timestamp 1666464484
transform 1 0 2352 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_25
timestamp 1666464484
transform 1 0 4144 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_33
timestamp 1666464484
transform 1 0 5040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_37
timestamp 1666464484
transform 1 0 5488 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_53
timestamp 1666464484
transform 1 0 7280 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_55
timestamp 1666464484
transform 1 0 7504 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_90
timestamp 1666464484
transform 1 0 11424 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_96
timestamp 1666464484
transform 1 0 12096 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_100
timestamp 1666464484
transform 1 0 12544 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_104
timestamp 1666464484
transform 1 0 12992 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_108
timestamp 1666464484
transform 1 0 13440 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_124
timestamp 1666464484
transform 1 0 15232 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_126
timestamp 1666464484
transform 1 0 15456 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_161
timestamp 1666464484
transform 1 0 19376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_167
timestamp 1666464484
transform 1 0 20048 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_171
timestamp 1666464484
transform 1 0 20496 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_175
timestamp 1666464484
transform 1 0 20944 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1666464484
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1666464484
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1666464484
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1666464484
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1666464484
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1666464484
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1666464484
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1666464484
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1666464484
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1666464484
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_456
timestamp 1666464484
transform 1 0 52416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1666464484
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_463
timestamp 1666464484
transform 1 0 53200 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_479
timestamp 1666464484
transform 1 0 54992 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_483
timestamp 1666464484
transform 1 0 55440 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_485
timestamp 1666464484
transform 1 0 55664 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_488
timestamp 1666464484
transform 1 0 56000 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_492
timestamp 1666464484
transform 1 0 56448 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_508
timestamp 1666464484
transform 1 0 58240 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_2
timestamp 1666464484
transform 1 0 1568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_6
timestamp 1666464484
transform 1 0 2016 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_21
timestamp 1666464484
transform 1 0 3696 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_25
timestamp 1666464484
transform 1 0 4144 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_33
timestamp 1666464484
transform 1 0 5040 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_37
timestamp 1666464484
transform 1 0 5488 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_52
timestamp 1666464484
transform 1 0 7168 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_56
timestamp 1666464484
transform 1 0 7616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_60
timestamp 1666464484
transform 1 0 8064 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_65
timestamp 1666464484
transform 1 0 8624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1666464484
transform 1 0 9072 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_72
timestamp 1666464484
transform 1 0 9408 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_80
timestamp 1666464484
transform 1 0 10304 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_84
timestamp 1666464484
transform 1 0 10752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_99
timestamp 1666464484
transform 1 0 12432 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_103
timestamp 1666464484
transform 1 0 12880 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_107
timestamp 1666464484
transform 1 0 13328 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1666464484
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_142
timestamp 1666464484
transform 1 0 17248 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_157
timestamp 1666464484
transform 1 0 18928 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_161
timestamp 1666464484
transform 1 0 19376 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_169
timestamp 1666464484
transform 1 0 20272 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_173
timestamp 1666464484
transform 1 0 20720 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_177
timestamp 1666464484
transform 1 0 21168 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_185
timestamp 1666464484
transform 1 0 22064 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_191
timestamp 1666464484
transform 1 0 22736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_207
timestamp 1666464484
transform 1 0 24528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1666464484
transform 1 0 24752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1666464484
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_215
timestamp 1666464484
transform 1 0 25424 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_231
timestamp 1666464484
transform 1 0 27216 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_239
timestamp 1666464484
transform 1 0 28112 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_241
timestamp 1666464484
transform 1 0 28336 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_244
timestamp 1666464484
transform 1 0 28672 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_247
timestamp 1666464484
transform 1 0 29008 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_262
timestamp 1666464484
transform 1 0 30688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_266
timestamp 1666464484
transform 1 0 31136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_269
timestamp 1666464484
transform 1 0 31472 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_277
timestamp 1666464484
transform 1 0 32368 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_279
timestamp 1666464484
transform 1 0 32592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_282
timestamp 1666464484
transform 1 0 32928 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_290
timestamp 1666464484
transform 1 0 33824 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_294
timestamp 1666464484
transform 1 0 34272 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_296
timestamp 1666464484
transform 1 0 34496 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_299
timestamp 1666464484
transform 1 0 34832 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_307
timestamp 1666464484
transform 1 0 35728 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_317
timestamp 1666464484
transform 1 0 36848 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_323
timestamp 1666464484
transform 1 0 37520 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_331
timestamp 1666464484
transform 1 0 38416 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_349
timestamp 1666464484
transform 1 0 40432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_352
timestamp 1666464484
transform 1 0 40768 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1666464484
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_369
timestamp 1666464484
transform 1 0 42672 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_387
timestamp 1666464484
transform 1 0 44688 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_395
timestamp 1666464484
transform 1 0 45584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_401
timestamp 1666464484
transform 1 0 46256 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_409
timestamp 1666464484
transform 1 0 47152 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_417
timestamp 1666464484
transform 1 0 48048 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_419
timestamp 1666464484
transform 1 0 48272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_422
timestamp 1666464484
transform 1 0 48608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_426
timestamp 1666464484
transform 1 0 49056 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_428
timestamp 1666464484
transform 1 0 49280 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_431
timestamp 1666464484
transform 1 0 49616 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_447
timestamp 1666464484
transform 1 0 51408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_451
timestamp 1666464484
transform 1 0 51856 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_454
timestamp 1666464484
transform 1 0 52192 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_457
timestamp 1666464484
transform 1 0 52528 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_464
timestamp 1666464484
transform 1 0 53312 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_472
timestamp 1666464484
transform 1 0 54208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_476
timestamp 1666464484
transform 1 0 54656 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_478
timestamp 1666464484
transform 1 0 54880 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_481
timestamp 1666464484
transform 1 0 55216 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_489
timestamp 1666464484
transform 1 0 56112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_492
timestamp 1666464484
transform 1 0 56448 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_508
timestamp 1666464484
transform 1 0 58240 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1666464484
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1666464484
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1666464484
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1666464484
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1666464484
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1666464484
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1666464484
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1666464484
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1666464484
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1666464484
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1666464484
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1666464484
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1666464484
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1666464484
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1666464484
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1666464484
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1666464484
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1666464484
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1666464484
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1666464484
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1666464484
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1666464484
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1666464484
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1666464484
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1666464484
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1666464484
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1666464484
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1666464484
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1666464484
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1666464484
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1666464484
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1666464484
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1666464484
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1666464484
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1666464484
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1666464484
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1666464484
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1666464484
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1666464484
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1666464484
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1666464484
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1666464484
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1666464484
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1666464484
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1666464484
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1666464484
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1666464484
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1666464484
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1666464484
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1666464484
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1666464484
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1666464484
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1666464484
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1666464484
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1666464484
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1666464484
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1666464484
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1666464484
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1666464484
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1666464484
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1666464484
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1666464484
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1666464484
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1666464484
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1666464484
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1666464484
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1666464484
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1666464484
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1666464484
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1666464484
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1666464484
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1666464484
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1666464484
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1666464484
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1666464484
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1666464484
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1666464484
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1666464484
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1666464484
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1666464484
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1666464484
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1666464484
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1666464484
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1666464484
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1666464484
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1666464484
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1666464484
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1666464484
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1666464484
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1666464484
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1666464484
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1666464484
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1666464484
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1666464484
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1666464484
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1666464484
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1666464484
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1666464484
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1666464484
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1666464484
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1666464484
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1666464484
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1666464484
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1666464484
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1666464484
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1666464484
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1666464484
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1666464484
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1666464484
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1666464484
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1666464484
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1666464484
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1666464484
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1666464484
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1666464484
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1666464484
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1666464484
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1666464484
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1666464484
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1666464484
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1666464484
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1666464484
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1666464484
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1666464484
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1666464484
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1666464484
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1666464484
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1666464484
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1666464484
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1666464484
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1666464484
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1666464484
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1666464484
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1666464484
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1666464484
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1666464484
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1666464484
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1666464484
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1666464484
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1666464484
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1666464484
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1666464484
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1666464484
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1666464484
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1666464484
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1666464484
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1666464484
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1666464484
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1666464484
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1666464484
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1666464484
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1666464484
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1666464484
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1666464484
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1666464484
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1666464484
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1666464484
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1666464484
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1666464484
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1666464484
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1666464484
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1666464484
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1666464484
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1666464484
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1666464484
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1666464484
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1666464484
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1666464484
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1666464484
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1666464484
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1666464484
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1666464484
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1666464484
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1666464484
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1666464484
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1666464484
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1666464484
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1666464484
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1666464484
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1666464484
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1666464484
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1666464484
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1666464484
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1666464484
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1666464484
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1666464484
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1666464484
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1666464484
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1666464484
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1666464484
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1666464484
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1666464484
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1666464484
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1666464484
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1666464484
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1666464484
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1666464484
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1666464484
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1666464484
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1666464484
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1666464484
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1666464484
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1666464484
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1666464484
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1666464484
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1666464484
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1666464484
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1666464484
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1666464484
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1666464484
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1666464484
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1666464484
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1666464484
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1666464484
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1666464484
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1666464484
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1666464484
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1666464484
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1666464484
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1666464484
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1666464484
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1666464484
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1666464484
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1666464484
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1666464484
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1666464484
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1666464484
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1666464484
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1666464484
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1666464484
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1666464484
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1666464484
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1666464484
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1666464484
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1666464484
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1666464484
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1666464484
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1666464484
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1666464484
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1666464484
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1666464484
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1666464484
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1666464484
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1666464484
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1666464484
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1666464484
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1666464484
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1666464484
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1666464484
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1666464484
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1666464484
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1666464484
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _253_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 19152 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _254_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 17024 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _255_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 22512 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _256_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 42224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _257_
timestamp 1666464484
transform -1 0 37520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _258_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 34272 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _259_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 38976 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _260_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 35616 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _261_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 23968 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _262_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 25424 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _263_
timestamp 1666464484
transform 1 0 33712 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _264_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 48832 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _265_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 47712 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _266_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 48384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _267_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 39648 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _268_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 40992 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _269_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 54656 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _270_
timestamp 1666464484
transform -1 0 51968 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _271_
timestamp 1666464484
transform 1 0 38752 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _272_
timestamp 1666464484
transform -1 0 45808 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _273_
timestamp 1666464484
transform -1 0 42560 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _274_
timestamp 1666464484
transform 1 0 12096 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _275_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 14672 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _276_
timestamp 1666464484
transform -1 0 13888 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _277_
timestamp 1666464484
transform -1 0 12096 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _278_
timestamp 1666464484
transform 1 0 5040 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _279_
timestamp 1666464484
transform 1 0 9072 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _280_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 11536 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _281_
timestamp 1666464484
transform 1 0 32368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _282_
timestamp 1666464484
transform 1 0 30912 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _283_
timestamp 1666464484
transform 1 0 33488 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _284_
timestamp 1666464484
transform 1 0 34608 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _285_
timestamp 1666464484
transform -1 0 40432 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _286_
timestamp 1666464484
transform -1 0 37744 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _287_
timestamp 1666464484
transform 1 0 27216 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _288_
timestamp 1666464484
transform -1 0 44240 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _289_
timestamp 1666464484
transform -1 0 40656 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _290_
timestamp 1666464484
transform -1 0 40208 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _291_
timestamp 1666464484
transform -1 0 38752 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _292_
timestamp 1666464484
transform 1 0 18032 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _293_
timestamp 1666464484
transform -1 0 23296 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _294_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 50624 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _295_
timestamp 1666464484
transform -1 0 45808 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _296_
timestamp 1666464484
transform 1 0 35392 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _297_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 38864 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _298_
timestamp 1666464484
transform 1 0 25312 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _299_
timestamp 1666464484
transform -1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _300_
timestamp 1666464484
transform 1 0 29456 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _301_
timestamp 1666464484
transform 1 0 31696 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1666464484
transform 1 0 39424 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _303_
timestamp 1666464484
transform 1 0 8176 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _304_
timestamp 1666464484
transform 1 0 18928 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _305_
timestamp 1666464484
transform 1 0 34832 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _306_
timestamp 1666464484
transform -1 0 40656 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _307_
timestamp 1666464484
transform -1 0 24080 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _308_
timestamp 1666464484
transform 1 0 15344 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _309_
timestamp 1666464484
transform 1 0 24640 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _310_
timestamp 1666464484
transform -1 0 14896 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _311_
timestamp 1666464484
transform -1 0 13104 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _312_
timestamp 1666464484
transform 1 0 3584 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _313_
timestamp 1666464484
transform 1 0 12432 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _314_
timestamp 1666464484
transform 1 0 17584 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _315_
timestamp 1666464484
transform -1 0 20384 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _316_
timestamp 1666464484
transform 1 0 16464 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _317_
timestamp 1666464484
transform 1 0 17360 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _318_
timestamp 1666464484
transform 1 0 18928 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _319_
timestamp 1666464484
transform -1 0 37520 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _320_
timestamp 1666464484
transform -1 0 20048 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _321_
timestamp 1666464484
transform -1 0 17136 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _322_
timestamp 1666464484
transform -1 0 14112 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _323_
timestamp 1666464484
transform 1 0 14784 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _324_
timestamp 1666464484
transform 1 0 15792 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _325_
timestamp 1666464484
transform 1 0 35728 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _326_
timestamp 1666464484
transform -1 0 17136 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _327_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 12768 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _328_
timestamp 1666464484
transform 1 0 11984 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _329_
timestamp 1666464484
transform 1 0 3584 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _330_
timestamp 1666464484
transform -1 0 14448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _331_
timestamp 1666464484
transform 1 0 11760 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _332_
timestamp 1666464484
transform -1 0 22624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _333_
timestamp 1666464484
transform -1 0 29008 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _334_
timestamp 1666464484
transform -1 0 28896 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _335_
timestamp 1666464484
transform -1 0 28224 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _336_
timestamp 1666464484
transform 1 0 26880 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _337_
timestamp 1666464484
transform -1 0 31024 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _338_
timestamp 1666464484
transform -1 0 28000 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _339_
timestamp 1666464484
transform -1 0 28336 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _340_
timestamp 1666464484
transform 1 0 25536 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _341_
timestamp 1666464484
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _342_
timestamp 1666464484
transform -1 0 34160 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _343_
timestamp 1666464484
transform 1 0 32368 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _344_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 38976 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _345_
timestamp 1666464484
transform -1 0 42336 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _346_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 36176 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _347_
timestamp 1666464484
transform -1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _348_
timestamp 1666464484
transform -1 0 32816 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _349_
timestamp 1666464484
transform 1 0 35056 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _350_
timestamp 1666464484
transform 1 0 36064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _351_
timestamp 1666464484
transform -1 0 40320 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _352_
timestamp 1666464484
transform -1 0 40656 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _353_
timestamp 1666464484
transform 1 0 16576 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _354_
timestamp 1666464484
transform 1 0 19712 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _355_
timestamp 1666464484
transform -1 0 29008 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _356_
timestamp 1666464484
transform -1 0 21952 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _357_
timestamp 1666464484
transform -1 0 50288 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _358_
timestamp 1666464484
transform 1 0 22176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _359_
timestamp 1666464484
transform 1 0 3584 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _360_
timestamp 1666464484
transform 1 0 19152 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _361_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 23520 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _362_
timestamp 1666464484
transform 1 0 23072 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _363_
timestamp 1666464484
transform 1 0 5600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _364_
timestamp 1666464484
transform 1 0 17584 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _365_
timestamp 1666464484
transform -1 0 34608 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _366_
timestamp 1666464484
transform 1 0 33488 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _367_
timestamp 1666464484
transform -1 0 41440 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1666464484
transform -1 0 40880 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _369_
timestamp 1666464484
transform 1 0 42000 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _370_
timestamp 1666464484
transform -1 0 42672 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _371_
timestamp 1666464484
transform -1 0 41776 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _372_
timestamp 1666464484
transform -1 0 32480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _373_
timestamp 1666464484
transform -1 0 33600 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _374_
timestamp 1666464484
transform -1 0 31696 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _375_
timestamp 1666464484
transform -1 0 30912 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _376_
timestamp 1666464484
transform -1 0 38640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _377_
timestamp 1666464484
transform -1 0 31472 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _378_
timestamp 1666464484
transform -1 0 33936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _379_
timestamp 1666464484
transform 1 0 35504 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _380_
timestamp 1666464484
transform -1 0 33936 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _381_
timestamp 1666464484
transform -1 0 32032 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _382_
timestamp 1666464484
transform -1 0 28448 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _383_
timestamp 1666464484
transform 1 0 29120 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _384_
timestamp 1666464484
transform 1 0 34272 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _385_
timestamp 1666464484
transform 1 0 34496 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _386_
timestamp 1666464484
transform -1 0 39648 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _387_
timestamp 1666464484
transform -1 0 38752 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _388_
timestamp 1666464484
transform 1 0 42112 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _389_
timestamp 1666464484
transform 1 0 47152 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _390_
timestamp 1666464484
transform -1 0 50736 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _391_
timestamp 1666464484
transform -1 0 49728 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _392_
timestamp 1666464484
transform -1 0 46256 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _393_
timestamp 1666464484
transform -1 0 46928 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _394_
timestamp 1666464484
transform 1 0 47376 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _395_
timestamp 1666464484
transform 1 0 48272 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _396_
timestamp 1666464484
transform -1 0 46368 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _397_
timestamp 1666464484
transform -1 0 46368 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _398_
timestamp 1666464484
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _399_
timestamp 1666464484
transform 1 0 40320 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _400_
timestamp 1666464484
transform 1 0 41664 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _401_
timestamp 1666464484
transform 1 0 42560 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _402_
timestamp 1666464484
transform -1 0 44688 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _403_
timestamp 1666464484
transform -1 0 44016 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _404_
timestamp 1666464484
transform 1 0 33600 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _405_
timestamp 1666464484
transform 1 0 34608 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _406_
timestamp 1666464484
transform 1 0 38080 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _407_
timestamp 1666464484
transform 1 0 32144 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _408_
timestamp 1666464484
transform -1 0 36848 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _409_
timestamp 1666464484
transform -1 0 23744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _410_
timestamp 1666464484
transform 1 0 24080 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _411_
timestamp 1666464484
transform 1 0 29456 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _412_
timestamp 1666464484
transform 1 0 37632 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _413_
timestamp 1666464484
transform -1 0 39872 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _414_
timestamp 1666464484
transform -1 0 22624 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _415_
timestamp 1666464484
transform -1 0 29904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1666464484
transform 1 0 23856 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _417_
timestamp 1666464484
transform -1 0 27328 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _418_
timestamp 1666464484
transform -1 0 26768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _419_
timestamp 1666464484
transform -1 0 43792 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _420_
timestamp 1666464484
transform -1 0 25872 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _421_
timestamp 1666464484
transform -1 0 18480 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _422_
timestamp 1666464484
transform 1 0 19488 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _423_
timestamp 1666464484
transform 1 0 22848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _424_
timestamp 1666464484
transform 1 0 28448 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _425_
timestamp 1666464484
transform 1 0 22288 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _426_
timestamp 1666464484
transform -1 0 25536 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _427_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 41888 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _428_
timestamp 1666464484
transform -1 0 36288 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _429_
timestamp 1666464484
transform -1 0 28224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _430_
timestamp 1666464484
transform -1 0 28896 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _431_
timestamp 1666464484
transform -1 0 31696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _432_
timestamp 1666464484
transform -1 0 27664 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _433_
timestamp 1666464484
transform -1 0 30688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _434_
timestamp 1666464484
transform -1 0 28000 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _435_
timestamp 1666464484
transform -1 0 27888 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _436_
timestamp 1666464484
transform -1 0 29680 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _437_
timestamp 1666464484
transform -1 0 28896 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _438_
timestamp 1666464484
transform -1 0 29008 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _439_
timestamp 1666464484
transform -1 0 36624 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _440_
timestamp 1666464484
transform -1 0 27552 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _441_
timestamp 1666464484
transform -1 0 30016 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _442_
timestamp 1666464484
transform -1 0 30464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _443_
timestamp 1666464484
transform -1 0 28784 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _444_
timestamp 1666464484
transform -1 0 30912 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _445_
timestamp 1666464484
transform -1 0 27552 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _446_
timestamp 1666464484
transform -1 0 32816 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _447_
timestamp 1666464484
transform -1 0 32368 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _448_
timestamp 1666464484
transform -1 0 32144 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _449_
timestamp 1666464484
transform -1 0 32144 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _450_
timestamp 1666464484
transform -1 0 36624 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _451_
timestamp 1666464484
transform -1 0 29344 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _452_
timestamp 1666464484
transform -1 0 30576 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _453_
timestamp 1666464484
transform -1 0 28672 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _454_
timestamp 1666464484
transform -1 0 31248 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _455_
timestamp 1666464484
transform -1 0 31696 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _456_
timestamp 1666464484
transform -1 0 31360 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _457_
timestamp 1666464484
transform -1 0 31696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _458_
timestamp 1666464484
transform -1 0 31360 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _459_
timestamp 1666464484
transform -1 0 32368 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _460_
timestamp 1666464484
transform -1 0 31808 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _461_
timestamp 1666464484
transform -1 0 34608 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _462_
timestamp 1666464484
transform -1 0 34272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _463_
timestamp 1666464484
transform -1 0 50288 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _464_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 9856 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _465_
timestamp 1666464484
transform -1 0 10976 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _466_
timestamp 1666464484
transform -1 0 10192 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _467_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 3584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _468_
timestamp 1666464484
transform 1 0 4480 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _469_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 9632 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _470_
timestamp 1666464484
transform 1 0 11536 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _471_
timestamp 1666464484
transform 1 0 41104 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _472_
timestamp 1666464484
transform 1 0 39424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _473_
timestamp 1666464484
transform 1 0 3584 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _474_
timestamp 1666464484
transform 1 0 3696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _475_
timestamp 1666464484
transform 1 0 7168 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _476_
timestamp 1666464484
transform 1 0 50736 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _477_
timestamp 1666464484
transform -1 0 12208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _478_
timestamp 1666464484
transform -1 0 11536 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _479_
timestamp 1666464484
transform 1 0 10416 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _480_
timestamp 1666464484
transform 1 0 11200 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _481_
timestamp 1666464484
transform -1 0 6496 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _482_
timestamp 1666464484
transform -1 0 11536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _483_
timestamp 1666464484
transform 1 0 9968 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _484_
timestamp 1666464484
transform 1 0 9408 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _485_
timestamp 1666464484
transform -1 0 12320 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1666464484
transform -1 0 11760 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _487_
timestamp 1666464484
transform -1 0 11312 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _488_
timestamp 1666464484
transform -1 0 35280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _489_
timestamp 1666464484
transform -1 0 10976 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _490_
timestamp 1666464484
transform 1 0 7840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _491_
timestamp 1666464484
transform -1 0 12208 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _492_
timestamp 1666464484
transform 1 0 8624 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _493_
timestamp 1666464484
transform 1 0 10080 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _494_
timestamp 1666464484
transform 1 0 4592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _495_
timestamp 1666464484
transform 1 0 9632 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _496_
timestamp 1666464484
transform -1 0 9408 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _497_
timestamp 1666464484
transform -1 0 4256 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _498_
timestamp 1666464484
transform 1 0 3696 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _499_
timestamp 1666464484
transform -1 0 38192 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _500_
timestamp 1666464484
transform -1 0 25984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _501_
timestamp 1666464484
transform -1 0 27216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _502_
timestamp 1666464484
transform -1 0 15344 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _503_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 26992 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _504_
timestamp 1666464484
transform 1 0 16240 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _505_
timestamp 1666464484
transform -1 0 19936 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _506_ GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 20384 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _507_
timestamp 1666464484
transform 1 0 20160 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _508_
timestamp 1666464484
transform -1 0 10752 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _509_
timestamp 1666464484
transform 1 0 20048 0 -1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _510_
timestamp 1666464484
transform -1 0 10976 0 1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _511_
timestamp 1666464484
transform 1 0 19040 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _512_
timestamp 1666464484
transform 1 0 16352 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _513_
timestamp 1666464484
transform -1 0 19936 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _514_
timestamp 1666464484
transform 1 0 20272 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _515_
timestamp 1666464484
transform -1 0 11424 0 1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _516_
timestamp 1666464484
transform 1 0 20048 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _517_
timestamp 1666464484
transform 1 0 8400 0 1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _518_
timestamp 1666464484
transform 1 0 16240 0 1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _519_
timestamp 1666464484
transform 1 0 13552 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _520_
timestamp 1666464484
transform -1 0 11200 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _521_
timestamp 1666464484
transform 1 0 18928 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _522_
timestamp 1666464484
transform 1 0 14224 0 1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _523_
timestamp 1666464484
transform -1 0 9184 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _524_
timestamp 1666464484
transform -1 0 10416 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _525_
timestamp 1666464484
transform -1 0 10416 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _526_
timestamp 1666464484
transform 1 0 20384 0 -1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _527_
timestamp 1666464484
transform 1 0 15568 0 1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _528_
timestamp 1666464484
transform 1 0 19488 0 -1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _529_
timestamp 1666464484
transform -1 0 17136 0 -1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _530_
timestamp 1666464484
transform 1 0 8288 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _531_
timestamp 1666464484
transform 1 0 14896 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _532_
timestamp 1666464484
transform -1 0 9184 0 -1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _533_
timestamp 1666464484
transform 1 0 12992 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _534_
timestamp 1666464484
transform 1 0 7952 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _535_
timestamp 1666464484
transform -1 0 9184 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _536_
timestamp 1666464484
transform 1 0 6384 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _537_
timestamp 1666464484
transform 1 0 14784 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 13552 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1666464484
transform -1 0 15232 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1666464484
transform 1 0 15232 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1666464484
transform -1 0 15232 0 -1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1666464484
transform -1 0 20832 0 1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_69 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_70
timestamp 1666464484
transform 1 0 57792 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_71
timestamp 1666464484
transform 1 0 57792 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_72
timestamp 1666464484
transform -1 0 8624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_73
timestamp 1666464484
transform 1 0 57792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cntr_example_74
timestamp 1666464484
transform -1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1680 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform -1 0 58240 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform -1 0 58240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1666464484
transform -1 0 58240 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1666464484
transform -1 0 32368 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1666464484
transform -1 0 49392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1666464484
transform -1 0 58240 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1666464484
transform 1 0 1680 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1666464484
transform 1 0 1680 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1666464484
transform -1 0 58240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1666464484
transform -1 0 51184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1666464484
transform 1 0 1680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1666464484
transform -1 0 58240 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1666464484
transform 1 0 1680 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1666464484
transform 1 0 35056 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1666464484
transform -1 0 47152 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1666464484
transform 1 0 1680 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1666464484
transform 1 0 23632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1666464484
transform 1 0 1680 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1666464484
transform -1 0 58240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1666464484
transform -1 0 58240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1666464484
transform 1 0 1680 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1666464484
transform -1 0 58240 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1666464484
transform 1 0 19600 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1666464484
transform 1 0 37744 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1666464484
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1666464484
transform 1 0 1680 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1666464484
transform 1 0 21280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1666464484
transform -1 0 56112 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1666464484
transform -1 0 58240 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1666464484
transform 1 0 29680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1666464484
transform -1 0 53312 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1666464484
transform 1 0 41776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1666464484
transform 1 0 1680 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1666464484
transform 1 0 1680 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input36
timestamp 1666464484
transform -1 0 58240 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output37 GF180PDK/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 16464 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output38
timestamp 1666464484
transform -1 0 46368 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output39
timestamp 1666464484
transform 1 0 56672 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output40
timestamp 1666464484
transform -1 0 3248 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output41
timestamp 1666464484
transform 1 0 34944 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output42
timestamp 1666464484
transform -1 0 3696 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output43
timestamp 1666464484
transform 1 0 56560 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output44
timestamp 1666464484
transform -1 0 24528 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output45
timestamp 1666464484
transform 1 0 56672 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output46
timestamp 1666464484
transform 1 0 56672 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output47
timestamp 1666464484
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output48
timestamp 1666464484
transform -1 0 3248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output49
timestamp 1666464484
transform -1 0 18928 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output50
timestamp 1666464484
transform 1 0 29120 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output51
timestamp 1666464484
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output52
timestamp 1666464484
transform -1 0 3248 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output53
timestamp 1666464484
transform -1 0 3248 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output54
timestamp 1666464484
transform -1 0 27216 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output55
timestamp 1666464484
transform 1 0 41104 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output56
timestamp 1666464484
transform 1 0 56672 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output57
timestamp 1666464484
transform -1 0 12432 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output58
timestamp 1666464484
transform -1 0 11088 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output59
timestamp 1666464484
transform -1 0 4368 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output60
timestamp 1666464484
transform 1 0 56672 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output61
timestamp 1666464484
transform -1 0 3248 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output62
timestamp 1666464484
transform 1 0 17584 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output63
timestamp 1666464484
transform -1 0 3248 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output64
timestamp 1666464484
transform 1 0 56672 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output65
timestamp 1666464484
transform 1 0 33040 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output66
timestamp 1666464484
transform -1 0 3248 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output67
timestamp 1666464484
transform 1 0 49840 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output68
timestamp 1666464484
transform -1 0 7168 0 -1 56448
box -86 -86 1654 870
<< labels >>
flabel metal3 s 200 38248 800 38472 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 59200 20104 59800 20328 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 59200 22792 59800 23016 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 59200 8008 59800 8232 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 31528 59200 31752 59800 0 FreeSans 896 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 47656 200 47880 800 0 FreeSans 896 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal3 s 59200 37576 59800 37800 0 FreeSans 896 0 0 0 io_in[15]
port 6 nsew signal input
flabel metal3 s 200 29512 800 29736 0 FreeSans 896 0 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 200 41608 800 41832 0 FreeSans 896 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal3 s 59200 1960 59800 2184 0 FreeSans 896 0 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 50344 200 50568 800 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 200 35560 800 35784 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 59080 200 59304 800 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 200 56392 800 56616 0 FreeSans 896 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34888 59200 35112 59800 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 46312 59200 46536 59800 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 200 44296 800 44520 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 23464 200 23688 800 0 FreeSans 896 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 200 8680 800 8904 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 59200 16744 59800 16968 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 59200 40936 59800 41160 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 200 14728 800 14952 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 59200 49672 59800 49896 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 19432 59200 19656 59800 0 FreeSans 896 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 37576 59200 37800 59800 0 FreeSans 896 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 200 59080 800 59304 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 38248 200 38472 800 0 FreeSans 896 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 59200 46984 59800 47208 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 59200 52360 59800 52584 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53704 200 53928 800 0 FreeSans 896 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 43624 59200 43848 59800 0 FreeSans 896 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 5320 200 5544 800 0 FreeSans 896 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 200 50344 800 50568 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 20776 200 21000 800 0 FreeSans 896 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 55720 59200 55944 59800 0 FreeSans 896 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 59200 43624 59800 43848 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 29512 200 29736 800 0 FreeSans 896 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 52360 59200 52584 59800 0 FreeSans 896 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 14728 200 14952 800 0 FreeSans 896 90 0 0 io_out[0]
port 38 nsew signal tristate
flabel metal2 s 44296 200 44520 800 0 FreeSans 896 90 0 0 io_out[10]
port 39 nsew signal tristate
flabel metal3 s 59200 14056 59800 14280 0 FreeSans 896 0 0 0 io_out[11]
port 40 nsew signal tristate
flabel metal3 s 200 47656 800 47880 0 FreeSans 896 0 0 0 io_out[12]
port 41 nsew signal tristate
flabel metal2 s 35560 200 35784 800 0 FreeSans 896 90 0 0 io_out[13]
port 42 nsew signal tristate
flabel metal2 s 1960 59200 2184 59800 0 FreeSans 896 90 0 0 io_out[14]
port 43 nsew signal tristate
flabel metal2 s 56392 200 56616 800 0 FreeSans 896 90 0 0 io_out[15]
port 44 nsew signal tristate
flabel metal2 s 22792 59200 23016 59800 0 FreeSans 896 90 0 0 io_out[16]
port 45 nsew signal tristate
flabel metal3 s 59200 10696 59800 10920 0 FreeSans 896 0 0 0 io_out[17]
port 46 nsew signal tristate
flabel metal3 s 59200 25480 59800 25704 0 FreeSans 896 0 0 0 io_out[18]
port 47 nsew signal tristate
flabel metal3 s 200 11368 800 11592 0 FreeSans 896 0 0 0 io_out[19]
port 48 nsew signal tristate
flabel metal3 s 200 2632 800 2856 0 FreeSans 896 0 0 0 io_out[1]
port 49 nsew signal tristate
flabel metal2 s 16744 59200 16968 59800 0 FreeSans 896 90 0 0 io_out[20]
port 50 nsew signal tristate
flabel metal2 s 28840 59200 29064 59800 0 FreeSans 896 90 0 0 io_out[21]
port 51 nsew signal tristate
flabel metal3 s 200 5320 800 5544 0 FreeSans 896 0 0 0 io_out[22]
port 52 nsew signal tristate
flabel metal2 s -56 200 168 800 0 FreeSans 896 90 0 0 io_out[23]
port 53 nsew signal tristate
flabel metal3 s 200 32200 800 32424 0 FreeSans 896 0 0 0 io_out[24]
port 54 nsew signal tristate
flabel metal2 s 25480 59200 25704 59800 0 FreeSans 896 90 0 0 io_out[25]
port 55 nsew signal tristate
flabel metal2 s 40936 59200 41160 59800 0 FreeSans 896 90 0 0 io_out[26]
port 56 nsew signal tristate
flabel metal2 s 58408 59200 58632 59800 0 FreeSans 896 90 0 0 io_out[27]
port 57 nsew signal tristate
flabel metal2 s 10696 59200 10920 59800 0 FreeSans 896 90 0 0 io_out[28]
port 58 nsew signal tristate
flabel metal2 s 8680 200 8904 800 0 FreeSans 896 90 0 0 io_out[29]
port 59 nsew signal tristate
flabel metal2 s 2632 200 2856 800 0 FreeSans 896 90 0 0 io_out[2]
port 60 nsew signal tristate
flabel metal3 s 59200 58408 59800 58632 0 FreeSans 896 0 0 0 io_out[30]
port 61 nsew signal tristate
flabel metal3 s 200 23464 800 23688 0 FreeSans 896 0 0 0 io_out[31]
port 62 nsew signal tristate
flabel metal2 s 26824 200 27048 800 0 FreeSans 896 90 0 0 io_out[32]
port 63 nsew signal tristate
flabel metal3 s 59200 55720 59800 55944 0 FreeSans 896 0 0 0 io_out[33]
port 64 nsew signal tristate
flabel metal3 s 59200 4648 59800 4872 0 FreeSans 896 0 0 0 io_out[34]
port 65 nsew signal tristate
flabel metal2 s 8008 59200 8232 59800 0 FreeSans 896 90 0 0 io_out[35]
port 66 nsew signal tristate
flabel metal3 s 59200 31528 59800 31752 0 FreeSans 896 0 0 0 io_out[36]
port 67 nsew signal tristate
flabel metal2 s 11368 200 11592 800 0 FreeSans 896 90 0 0 io_out[37]
port 68 nsew signal tristate
flabel metal2 s 17416 200 17640 800 0 FreeSans 896 90 0 0 io_out[3]
port 69 nsew signal tristate
flabel metal3 s 200 26152 800 26376 0 FreeSans 896 0 0 0 io_out[4]
port 70 nsew signal tristate
flabel metal3 s 59200 34888 59800 35112 0 FreeSans 896 0 0 0 io_out[5]
port 71 nsew signal tristate
flabel metal2 s 32200 200 32424 800 0 FreeSans 896 90 0 0 io_out[6]
port 72 nsew signal tristate
flabel metal3 s 200 20776 800 21000 0 FreeSans 896 0 0 0 io_out[7]
port 73 nsew signal tristate
flabel metal2 s 49672 59200 49896 59800 0 FreeSans 896 90 0 0 io_out[8]
port 74 nsew signal tristate
flabel metal2 s 4648 59200 4872 59800 0 FreeSans 896 90 0 0 io_out[9]
port 75 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 76 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 76 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 77 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 77 nsew ground bidirectional
flabel metal2 s 14056 59200 14280 59800 0 FreeSans 896 90 0 0 wb_clk_i
port 78 nsew signal input
flabel metal2 s 41608 200 41832 800 0 FreeSans 896 90 0 0 wb_rst_i
port 79 nsew signal input
flabel metal3 s 200 17416 800 17640 0 FreeSans 896 0 0 0 wbs_cyc_i
port 80 nsew signal input
flabel metal3 s 200 53032 800 53256 0 FreeSans 896 0 0 0 wbs_stb_i
port 81 nsew signal input
flabel metal3 s 59200 28840 59800 29064 0 FreeSans 896 0 0 0 wbs_we_i
port 82 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 23464 47040 23464 47040 0 _000_
rlabel metal2 28616 47152 28616 47152 0 _001_
rlabel metal2 7784 45472 7784 45472 0 _002_
rlabel metal3 25312 53592 25312 53592 0 _003_
rlabel metal2 30408 52024 30408 52024 0 _004_
rlabel metal2 27720 43512 27720 43512 0 _005_
rlabel metal2 27552 47992 27552 47992 0 _006_
rlabel metal2 16968 46144 16968 46144 0 _007_
rlabel metal2 28616 46032 28616 46032 0 _008_
rlabel metal2 28728 53984 28728 53984 0 _009_
rlabel metal2 27272 44688 27272 44688 0 _010_
rlabel metal2 29736 53200 29736 53200 0 _011_
rlabel metal2 22176 52136 22176 52136 0 _012_
rlabel metal2 28504 43736 28504 43736 0 _013_
rlabel metal2 30576 45640 30576 45640 0 _014_
rlabel metal3 24696 50904 24696 50904 0 _015_
rlabel metal2 17416 53592 17416 53592 0 _016_
rlabel metal2 9800 44856 9800 44856 0 _017_
rlabel metal3 31864 40432 31864 40432 0 _018_
rlabel metal3 7924 48776 7924 48776 0 _019_
rlabel metal3 26264 53144 26264 53144 0 _020_
rlabel metal2 20888 54488 20888 54488 0 _021_
rlabel metal2 22680 51856 22680 51856 0 _022_
rlabel metal2 30968 53200 30968 53200 0 _023_
rlabel metal2 31416 49000 31416 49000 0 _024_
rlabel metal2 31080 52080 31080 52080 0 _025_
rlabel metal2 31416 52472 31416 52472 0 _026_
rlabel metal2 17752 43960 17752 43960 0 _027_
rlabel metal2 11144 49952 11144 49952 0 _028_
rlabel metal2 31528 43176 31528 43176 0 _029_
rlabel metal2 9576 43064 9576 43064 0 _030_
rlabel metal2 33992 44912 33992 44912 0 _031_
rlabel metal2 24584 46480 24584 46480 0 _032_
rlabel metal2 24416 44968 24416 44968 0 _033_
rlabel metal3 12824 45864 12824 45864 0 _034_
rlabel metal2 20776 54432 20776 54432 0 _035_
rlabel metal3 13552 52248 13552 52248 0 _036_
rlabel metal2 23240 39592 23240 39592 0 _037_
rlabel metal3 18760 39032 18760 39032 0 _038_
rlabel metal3 20048 45864 20048 45864 0 _039_
rlabel metal2 30072 44296 30072 44296 0 _040_
rlabel metal2 30408 47488 30408 47488 0 _041_
rlabel metal2 40824 38360 40824 38360 0 _042_
rlabel metal3 10808 53704 10808 53704 0 _043_
rlabel metal2 18984 51688 18984 51688 0 _044_
rlabel metal2 39704 36008 39704 36008 0 _045_
rlabel metal3 11368 44296 11368 44296 0 _046_
rlabel metal2 28392 46676 28392 46676 0 _047_
rlabel metal2 13832 51072 13832 51072 0 _048_
rlabel metal2 10808 43288 10808 43288 0 _049_
rlabel metal2 9800 41104 9800 41104 0 _050_
rlabel metal3 12096 48776 12096 48776 0 _051_
rlabel metal2 24584 52416 24584 52416 0 _052_
rlabel metal2 20328 54768 20328 54768 0 _053_
rlabel metal2 37800 47712 37800 47712 0 _054_
rlabel metal3 17360 52920 17360 52920 0 _055_
rlabel metal2 9072 47432 9072 47432 0 _056_
rlabel metal3 17696 50568 17696 50568 0 _057_
rlabel metal2 10304 52808 10304 52808 0 _058_
rlabel metal2 12712 43008 12712 43008 0 _059_
rlabel metal3 11984 50456 11984 50456 0 _060_
rlabel metal3 9912 45080 9912 45080 0 _061_
rlabel metal2 7112 42504 7112 42504 0 _062_
rlabel metal3 11256 44072 11256 44072 0 _063_
rlabel metal3 27552 26488 27552 26488 0 _064_
rlabel metal2 22064 23688 22064 23688 0 _065_
rlabel metal2 9912 23240 9912 23240 0 _066_
rlabel metal2 10584 35672 10584 35672 0 _067_
rlabel metal2 4312 23464 4312 23464 0 _068_
rlabel metal3 4088 51128 4088 51128 0 _069_
rlabel metal2 24696 26488 24696 26488 0 _070_
rlabel metal3 38136 50456 38136 50456 0 _071_
rlabel metal3 40040 31528 40040 31528 0 _072_
rlabel metal2 4368 53704 4368 53704 0 _073_
rlabel metal2 3696 53480 3696 53480 0 _074_
rlabel metal3 6104 38584 6104 38584 0 _075_
rlabel metal2 51576 51240 51576 51240 0 _076_
rlabel metal2 10920 25760 10920 25760 0 _077_
rlabel metal2 10640 25592 10640 25592 0 _078_
rlabel metal2 11536 25592 11536 25592 0 _079_
rlabel metal2 11480 27384 11480 27384 0 _080_
rlabel metal3 8120 27720 8120 27720 0 _081_
rlabel metal2 10920 26264 10920 26264 0 _082_
rlabel metal3 10136 32760 10136 32760 0 _083_
rlabel metal3 11256 32648 11256 32648 0 _084_
rlabel metal2 11256 30968 11256 30968 0 _085_
rlabel metal2 10752 29624 10752 29624 0 _086_
rlabel metal3 34440 40152 34440 40152 0 _087_
rlabel metal3 9296 34216 9296 34216 0 _088_
rlabel metal2 9016 36512 9016 36512 0 _089_
rlabel metal3 9688 34776 9688 34776 0 _090_
rlabel metal2 10024 34384 10024 34384 0 _091_
rlabel metal3 7392 33992 7392 33992 0 _092_
rlabel metal3 6496 36568 6496 36568 0 _093_
rlabel metal2 3752 45052 3752 45052 0 _094_
rlabel metal3 30968 45528 30968 45528 0 _095_
rlabel metal3 20384 37240 20384 37240 0 _096_
rlabel metal2 26712 36400 26712 36400 0 _097_
rlabel metal3 26264 37240 26264 37240 0 _098_
rlabel metal3 30856 40488 30856 40488 0 _099_
rlabel metal2 18760 28672 18760 28672 0 _100_
rlabel metal2 18984 29736 18984 29736 0 _101_
rlabel metal3 20664 28616 20664 28616 0 _102_
rlabel metal2 22344 23464 22344 23464 0 _103_
rlabel metal2 25144 25424 25144 25424 0 _104_
rlabel metal2 41888 35560 41888 35560 0 _105_
rlabel metal2 35168 33544 35168 33544 0 _106_
rlabel metal2 38808 38808 38808 38808 0 _107_
rlabel metal3 36064 36568 36064 36568 0 _108_
rlabel metal2 24248 28560 24248 28560 0 _109_
rlabel metal2 27944 40712 27944 40712 0 _110_
rlabel metal2 53144 51632 53144 51632 0 _111_
rlabel metal2 46648 48496 46648 48496 0 _112_
rlabel metal2 47992 46704 47992 46704 0 _113_
rlabel metal2 48104 46592 48104 46592 0 _114_
rlabel metal2 41608 48832 41608 48832 0 _115_
rlabel metal2 40824 51744 40824 51744 0 _116_
rlabel metal3 52640 52136 52640 52136 0 _117_
rlabel metal2 51464 52976 51464 52976 0 _118_
rlabel metal3 40824 53816 40824 53816 0 _119_
rlabel metal3 43624 53480 43624 53480 0 _120_
rlabel metal3 11144 30184 11144 30184 0 _121_
rlabel metal2 13048 31416 13048 31416 0 _122_
rlabel metal2 12712 31360 12712 31360 0 _123_
rlabel metal3 10640 30408 10640 30408 0 _124_
rlabel metal3 7392 30408 7392 30408 0 _125_
rlabel metal3 37576 45864 37576 45864 0 _126_
rlabel metal2 34216 43176 34216 43176 0 _127_
rlabel metal2 31416 41328 31416 41328 0 _128_
rlabel metal2 34720 42840 34720 42840 0 _129_
rlabel metal3 36232 43288 36232 43288 0 _130_
rlabel metal2 39928 40936 39928 40936 0 _131_
rlabel metal3 29344 41272 29344 41272 0 _132_
rlabel metal3 41776 50792 41776 50792 0 _133_
rlabel metal2 38360 46592 38360 46592 0 _134_
rlabel metal3 39256 45304 39256 45304 0 _135_
rlabel metal3 22176 33096 22176 33096 0 _136_
rlabel metal2 22176 23352 22176 23352 0 _137_
rlabel metal2 46088 36400 46088 36400 0 _138_
rlabel metal2 45528 40768 45528 40768 0 _139_
rlabel metal3 37744 38920 37744 38920 0 _140_
rlabel metal2 39256 36456 39256 36456 0 _141_
rlabel metal2 26488 36008 26488 36008 0 _142_
rlabel metal2 28840 39704 28840 39704 0 _143_
rlabel metal3 30800 40264 30800 40264 0 _144_
rlabel metal2 19320 37352 19320 37352 0 _145_
rlabel metal2 4536 48608 4536 48608 0 _146_
rlabel metal2 18984 37016 18984 37016 0 _147_
rlabel metal2 40208 34888 40208 34888 0 _148_
rlabel metal2 39928 34440 39928 34440 0 _149_
rlabel metal2 23688 33488 23688 33488 0 _150_
rlabel metal2 39592 36008 39592 36008 0 _151_
rlabel metal2 13720 37240 13720 37240 0 _152_
rlabel metal2 12824 37520 12824 37520 0 _153_
rlabel metal3 4536 49000 4536 49000 0 _154_
rlabel metal3 18536 36456 18536 36456 0 _155_
rlabel metal2 18088 30968 18088 30968 0 _156_
rlabel metal2 17192 32648 17192 32648 0 _157_
rlabel metal3 18816 34776 18816 34776 0 _158_
rlabel metal2 19544 35112 19544 35112 0 _159_
rlabel metal2 37184 40376 37184 40376 0 _160_
rlabel metal3 16576 35672 16576 35672 0 _161_
rlabel metal2 15176 33824 15176 33824 0 _162_
rlabel metal2 15960 35672 15960 35672 0 _163_
rlabel metal2 16744 35952 16744 35952 0 _164_
rlabel metal4 30968 45528 30968 45528 0 _165_
rlabel metal2 11984 28840 11984 28840 0 _166_
rlabel metal2 12208 32760 12208 32760 0 _167_
rlabel metal3 4368 47320 4368 47320 0 _168_
rlabel metal3 13384 35896 13384 35896 0 _169_
rlabel metal2 26040 27216 26040 27216 0 _170_
rlabel metal3 28000 27048 28000 27048 0 _171_
rlabel metal2 28504 28952 28504 28952 0 _172_
rlabel metal2 26992 26376 26992 26376 0 _173_
rlabel metal2 27440 26152 27440 26152 0 _174_
rlabel metal3 29344 31864 29344 31864 0 _175_
rlabel metal2 27496 32872 27496 32872 0 _176_
rlabel metal3 28952 44968 28952 44968 0 _177_
rlabel metal2 39368 28672 39368 28672 0 _178_
rlabel metal2 33768 27888 33768 27888 0 _179_
rlabel metal2 39144 28392 39144 28392 0 _180_
rlabel metal3 40768 26376 40768 26376 0 _181_
rlabel metal2 42056 26712 42056 26712 0 _182_
rlabel metal2 39816 35616 39816 35616 0 _183_
rlabel metal2 22680 32480 22680 32480 0 _184_
rlabel metal2 35560 32928 35560 32928 0 _185_
rlabel metal2 40264 35280 40264 35280 0 _186_
rlabel metal3 40208 31976 40208 31976 0 _187_
rlabel metal3 29232 45080 29232 45080 0 _188_
rlabel metal3 20832 33880 20832 33880 0 _189_
rlabel metal2 24696 27664 24696 27664 0 _190_
rlabel metal3 21840 32536 21840 32536 0 _191_
rlabel metal2 31024 39032 31024 39032 0 _192_
rlabel metal2 22568 33992 22568 33992 0 _193_
rlabel metal2 3976 43792 3976 43792 0 _194_
rlabel metal2 23240 28616 23240 28616 0 _195_
rlabel metal2 23352 28448 23352 28448 0 _196_
rlabel metal2 17080 29960 17080 29960 0 _197_
rlabel metal3 33824 36680 33824 36680 0 _198_
rlabel metal3 41440 38136 41440 38136 0 _199_
rlabel metal2 40712 37576 40712 37576 0 _200_
rlabel metal3 40992 36680 40992 36680 0 _201_
rlabel metal2 28224 53480 28224 53480 0 _202_
rlabel metal3 41888 36568 41888 36568 0 _203_
rlabel via2 31416 36456 31416 36456 0 _204_
rlabel metal3 32200 38024 32200 38024 0 _205_
rlabel metal2 31024 38024 31024 38024 0 _206_
rlabel metal2 31080 37240 31080 37240 0 _207_
rlabel metal2 31528 35504 31528 35504 0 _208_
rlabel metal3 30352 45304 30352 45304 0 _209_
rlabel metal2 33712 39704 33712 39704 0 _210_
rlabel metal2 31808 39592 31808 39592 0 _211_
rlabel metal2 31640 40768 31640 40768 0 _212_
rlabel metal2 27608 46424 27608 46424 0 _213_
rlabel metal2 34552 34608 34552 34608 0 _214_
rlabel metal3 36624 33544 36624 33544 0 _215_
rlabel metal3 38976 31864 38976 31864 0 _216_
rlabel metal2 47544 39984 47544 39984 0 _217_
rlabel metal3 49224 39480 49224 39480 0 _218_
rlabel metal2 49560 36904 49560 36904 0 _219_
rlabel metal3 47992 35672 47992 35672 0 _220_
rlabel metal2 45976 34384 45976 34384 0 _221_
rlabel metal2 48328 39704 48328 39704 0 _222_
rlabel metal3 47264 38808 47264 38808 0 _223_
rlabel metal2 46144 35000 46144 35000 0 _224_
rlabel metal2 40824 45360 40824 45360 0 _225_
rlabel metal3 41216 39816 41216 39816 0 _226_
rlabel metal2 42392 41160 42392 41160 0 _227_
rlabel metal3 43232 41272 43232 41272 0 _228_
rlabel metal2 43848 48104 43848 48104 0 _229_
rlabel metal2 34944 39480 34944 39480 0 _230_
rlabel metal3 36624 39592 36624 39592 0 _231_
rlabel metal3 37408 39704 37408 39704 0 _232_
rlabel metal2 34328 40320 34328 40320 0 _233_
rlabel metal2 23352 34608 23352 34608 0 _234_
rlabel metal2 24864 24920 24864 24920 0 _235_
rlabel metal3 33432 31752 33432 31752 0 _236_
rlabel metal2 38472 31752 38472 31752 0 _237_
rlabel metal4 39480 36400 39480 36400 0 _238_
rlabel metal2 25032 35672 25032 35672 0 _239_
rlabel metal2 24080 25704 24080 25704 0 _240_
rlabel metal2 26712 32872 26712 32872 0 _241_
rlabel metal2 26320 32760 26320 32760 0 _242_
rlabel metal2 43064 52696 43064 52696 0 _243_
rlabel metal2 18088 23968 18088 23968 0 _244_
rlabel metal2 19712 24920 19712 24920 0 _245_
rlabel metal3 24192 27048 24192 27048 0 _246_
rlabel metal2 25368 29064 25368 29064 0 _247_
rlabel metal3 23632 26936 23632 26936 0 _248_
rlabel metal2 41384 29344 41384 29344 0 _249_
rlabel metal2 27496 54096 27496 54096 0 _250_
rlabel metal2 27496 52136 27496 52136 0 _251_
rlabel metal3 29008 52248 29008 52248 0 _252_
rlabel metal2 15064 41888 15064 41888 0 clknet_0_wb_clk_i
rlabel metal2 8848 45080 8848 45080 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 15064 43988 15064 43988 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 8232 51744 8232 51744 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 20552 52584 20552 52584 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 1848 38192 1848 38192 0 io_in[0]
rlabel metal2 58072 20496 58072 20496 0 io_in[10]
rlabel metal2 58072 23072 58072 23072 0 io_in[11]
rlabel metal3 58674 8120 58674 8120 0 io_in[12]
rlabel metal2 31472 56280 31472 56280 0 io_in[13]
rlabel metal2 48216 2072 48216 2072 0 io_in[14]
rlabel metal2 58072 37856 58072 37856 0 io_in[15]
rlabel metal3 1302 29624 1302 29624 0 io_in[16]
rlabel metal2 1848 41888 1848 41888 0 io_in[17]
rlabel metal2 58072 3584 58072 3584 0 io_in[18]
rlabel metal2 50344 3416 50344 3416 0 io_in[19]
rlabel metal3 1246 35784 1246 35784 0 io_in[1]
rlabel metal2 58128 4984 58128 4984 0 io_in[20]
rlabel metal2 1848 54936 1848 54936 0 io_in[21]
rlabel metal2 34832 56280 34832 56280 0 io_in[22]
rlabel metal2 46256 56280 46256 56280 0 io_in[23]
rlabel metal3 1302 44408 1302 44408 0 io_in[24]
rlabel metal2 23464 3416 23464 3416 0 io_in[25]
rlabel metal3 1302 8680 1302 8680 0 io_in[26]
rlabel metal2 58072 17248 58072 17248 0 io_in[27]
rlabel metal3 58674 41048 58674 41048 0 io_in[28]
rlabel metal2 1848 14672 1848 14672 0 io_in[29]
rlabel metal3 58688 50456 58688 50456 0 io_in[2]
rlabel metal2 19376 56280 19376 56280 0 io_in[30]
rlabel metal2 37520 56280 37520 56280 0 io_in[31]
rlabel metal2 5208 3416 5208 3416 0 io_in[3]
rlabel metal3 1302 50456 1302 50456 0 io_in[4]
rlabel metal2 20776 2086 20776 2086 0 io_in[5]
rlabel metal2 55944 57722 55944 57722 0 io_in[6]
rlabel metal2 58072 44016 58072 44016 0 io_in[7]
rlabel metal2 29456 3416 29456 3416 0 io_in[8]
rlabel metal2 52248 56280 52248 56280 0 io_in[9]
rlabel metal2 14952 2198 14952 2198 0 io_out[0]
rlabel metal2 44520 798 44520 798 0 io_out[10]
rlabel metal2 57736 14336 57736 14336 0 io_out[11]
rlabel metal3 1414 47880 1414 47880 0 io_out[12]
rlabel metal2 35784 2198 35784 2198 0 io_out[13]
rlabel metal2 2632 57736 2632 57736 0 io_out[14]
rlabel metal2 56616 2086 56616 2086 0 io_out[15]
rlabel metal2 23464 57736 23464 57736 0 io_out[16]
rlabel metal2 57736 11088 57736 11088 0 io_out[17]
rlabel metal3 58562 25592 58562 25592 0 io_out[18]
rlabel metal3 1414 11592 1414 11592 0 io_out[19]
rlabel metal3 1414 2856 1414 2856 0 io_out[1]
rlabel metal2 17752 57624 17752 57624 0 io_out[20]
rlabel metal2 29960 56280 29960 56280 0 io_out[21]
rlabel metal3 1414 5544 1414 5544 0 io_out[22]
rlabel metal2 168 798 168 798 0 io_out[23]
rlabel metal3 1414 32424 1414 32424 0 io_out[24]
rlabel metal2 26152 57736 26152 57736 0 io_out[25]
rlabel metal3 41664 56168 41664 56168 0 io_out[26]
rlabel metal2 57736 57736 57736 57736 0 io_out[27]
rlabel metal2 11368 57736 11368 57736 0 io_out[28]
rlabel metal2 8904 2086 8904 2086 0 io_out[29]
rlabel metal2 2856 798 2856 798 0 io_out[2]
rlabel metal3 58576 57736 58576 57736 0 io_out[30]
rlabel metal3 1470 23688 1470 23688 0 io_out[31]
rlabel metal2 17640 798 17640 798 0 io_out[3]
rlabel metal3 1470 26376 1470 26376 0 io_out[4]
rlabel metal3 58562 35000 58562 35000 0 io_out[5]
rlabel metal2 32424 2086 32424 2086 0 io_out[6]
rlabel metal3 1414 21000 1414 21000 0 io_out[7]
rlabel metal3 50288 55944 50288 55944 0 io_out[8]
rlabel metal3 5488 56168 5488 56168 0 io_out[9]
rlabel metal3 2856 46536 2856 46536 0 net1
rlabel metal3 40880 30856 40880 30856 0 net10
rlabel metal3 46536 3304 46536 3304 0 net11
rlabel metal2 2184 35224 2184 35224 0 net12
rlabel metal2 57680 4984 57680 4984 0 net13
rlabel metal3 3024 53032 3024 53032 0 net14
rlabel metal2 35896 47488 35896 47488 0 net15
rlabel metal2 46536 50316 46536 50316 0 net16
rlabel metal2 2184 47040 2184 47040 0 net17
rlabel metal4 24360 28280 24360 28280 0 net18
rlabel metal3 5096 26600 5096 26600 0 net19
rlabel metal2 46592 34664 46592 34664 0 net2
rlabel metal3 40824 44968 40824 44968 0 net20
rlabel metal2 40264 40320 40264 40320 0 net21
rlabel metal2 2240 15512 2240 15512 0 net22
rlabel metal2 57680 50344 57680 50344 0 net23
rlabel metal2 20216 54880 20216 54880 0 net24
rlabel metal3 39032 56168 39032 56168 0 net25
rlabel metal2 6216 3304 6216 3304 0 net26
rlabel metal2 2128 50344 2128 50344 0 net27
rlabel metal3 24976 3304 24976 3304 0 net28
rlabel metal3 49616 52808 49616 52808 0 net29
rlabel metal2 46704 33992 46704 33992 0 net3
rlabel metal3 40992 38024 40992 38024 0 net30
rlabel metal3 30912 3304 30912 3304 0 net31
rlabel metal2 44520 49952 44520 49952 0 net32
rlabel metal2 42168 3304 42168 3304 0 net33
rlabel metal2 2184 18088 2184 18088 0 net34
rlabel metal3 3416 51464 3416 51464 0 net35
rlabel metal3 49448 46536 49448 46536 0 net36
rlabel metal2 16520 4928 16520 4928 0 net37
rlabel metal2 45808 3528 45808 3528 0 net38
rlabel metal2 51352 23268 51352 23268 0 net39
rlabel metal3 39928 31640 39928 31640 0 net4
rlabel metal2 3304 46424 3304 46424 0 net40
rlabel metal2 34944 3528 34944 3528 0 net41
rlabel metal2 7840 51352 7840 51352 0 net42
rlabel metal3 56392 3528 56392 3528 0 net43
rlabel metal2 21840 24920 21840 24920 0 net44
rlabel metal2 27888 24920 27888 24920 0 net45
rlabel metal2 28672 24920 28672 24920 0 net46
rlabel metal2 28392 24976 28392 24976 0 net47
rlabel metal2 3472 4536 3472 4536 0 net48
rlabel metal3 21728 55944 21728 55944 0 net49
rlabel metal2 28336 53032 28336 53032 0 net5
rlabel metal3 28952 55160 28952 55160 0 net50
rlabel metal3 4984 6104 4984 6104 0 net51
rlabel metal3 4928 5208 4928 5208 0 net52
rlabel metal2 6496 48776 6496 48776 0 net53
rlabel metal3 25032 52696 25032 52696 0 net54
rlabel metal2 28224 47320 28224 47320 0 net55
rlabel metal2 38024 48160 38024 48160 0 net56
rlabel metal2 13328 52696 13328 52696 0 net57
rlabel metal3 11760 4536 11760 4536 0 net58
rlabel metal2 4368 4536 4368 4536 0 net59
rlabel metal2 48888 3248 48888 3248 0 net6
rlabel metal3 53424 52248 53424 52248 0 net60
rlabel metal3 4760 24024 4760 24024 0 net61
rlabel metal3 14336 3640 14336 3640 0 net62
rlabel metal2 3080 26992 3080 26992 0 net63
rlabel metal3 23576 25592 23576 25592 0 net64
rlabel metal2 23240 24976 23240 24976 0 net65
rlabel metal2 3528 22736 3528 22736 0 net66
rlabel metal2 23912 54264 23912 54264 0 net67
rlabel metal2 7224 46032 7224 46032 0 net68
rlabel metal2 27048 2030 27048 2030 0 net69
rlabel metal2 43512 37016 43512 37016 0 net7
rlabel metal2 58072 55048 58072 55048 0 net70
rlabel metal2 58072 5600 58072 5600 0 net71
rlabel metal2 8288 56280 8288 56280 0 net72
rlabel metal3 58674 31528 58674 31528 0 net73
rlabel metal2 11592 2030 11592 2030 0 net74
rlabel metal2 2184 30184 2184 30184 0 net8
rlabel metal3 2912 47096 2912 47096 0 net9
rlabel metal2 14056 53354 14056 53354 0 wb_clk_i
rlabel metal2 41552 3416 41552 3416 0 wb_rst_i
rlabel metal3 1302 17528 1302 17528 0 wbs_cyc_i
rlabel metal3 1302 53144 1302 53144 0 wbs_stb_i
rlabel metal2 58184 28784 58184 28784 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
