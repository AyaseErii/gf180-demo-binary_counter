VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cntr_example
  CLASS BLOCK ;
  FOREIGN cntr_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.240 4.000 192.360 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 100.520 299.000 101.640 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 113.960 299.000 115.080 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 40.040 299.000 41.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.640 296.000 158.760 299.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 1.000 239.400 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 187.880 299.000 189.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.560 4.000 148.680 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.040 4.000 209.160 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 9.800 299.000 10.920 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.720 1.000 252.840 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 177.800 4.000 178.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.400 1.000 296.520 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 281.960 4.000 283.080 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 296.000 175.560 299.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 296.000 232.680 299.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.480 4.000 222.600 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.320 1.000 118.440 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.400 4.000 44.520 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 83.720 299.000 84.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 204.680 299.000 205.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.640 4.000 74.760 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 248.360 299.000 249.480 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 296.000 98.280 299.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.880 296.000 189.000 299.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 295.400 4.000 296.520 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 1.000 192.360 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 234.920 299.000 236.040 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 261.800 299.000 262.920 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 1.000 269.640 4.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 296.000 219.240 299.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 1.000 27.720 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 251.720 4.000 252.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 1.000 105.000 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 296.000 279.720 299.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 218.120 299.000 219.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.560 1.000 148.680 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.800 296.000 262.920 299.000 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 1.000 74.760 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.480 1.000 222.600 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 70.280 299.000 71.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.280 4.000 239.400 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 1.000 178.920 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 296.000 10.920 299.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.960 1.000 283.080 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 296.000 115.080 299.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 53.480 299.000 54.600 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 127.400 299.000 128.520 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 56.840 4.000 57.960 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.160 4.000 14.280 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.720 296.000 84.840 299.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 296.000 145.320 299.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.600 4.000 27.720 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 1.000 0.840 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.000 4.000 162.120 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.400 296.000 128.520 299.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.680 296.000 205.800 299.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.040 296.000 293.160 299.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 296.000 54.600 299.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.400 1.000 44.520 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 1.000 14.280 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 292.040 299.000 293.160 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 117.320 4.000 118.440 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 1.000 135.240 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 278.600 299.000 279.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 23.240 299.000 24.360 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 296.000 41.160 299.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 157.640 299.000 158.760 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 1.000 57.960 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.080 1.000 88.200 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 130.760 4.000 131.880 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.440 299.000 175.560 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.000 1.000 162.120 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 103.880 4.000 105.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 296.000 249.480 299.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.240 296.000 24.360 299.000 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 296.000 71.400 299.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 1.000 209.160 4.000 ;
    END
  END wb_rst_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 87.080 4.000 88.200 ;
    END
  END wbs_cyc_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 265.160 4.000 266.280 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 144.200 299.000 145.320 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 0.700 295.700 9.500 296.660 ;
        RECT 11.220 295.700 22.940 296.660 ;
        RECT 24.660 295.700 39.740 296.660 ;
        RECT 41.460 295.700 53.180 296.660 ;
        RECT 54.900 295.700 69.980 296.660 ;
        RECT 71.700 295.700 83.420 296.660 ;
        RECT 85.140 295.700 96.860 296.660 ;
        RECT 98.580 295.700 113.660 296.660 ;
        RECT 115.380 295.700 127.100 296.660 ;
        RECT 128.820 295.700 143.900 296.660 ;
        RECT 145.620 295.700 157.340 296.660 ;
        RECT 159.060 295.700 174.140 296.660 ;
        RECT 175.860 295.700 187.580 296.660 ;
        RECT 189.300 295.700 204.380 296.660 ;
        RECT 206.100 295.700 217.820 296.660 ;
        RECT 219.540 295.700 231.260 296.660 ;
        RECT 232.980 295.700 248.060 296.660 ;
        RECT 249.780 295.700 261.500 296.660 ;
        RECT 263.220 295.700 278.300 296.660 ;
        RECT 280.020 295.700 291.740 296.660 ;
        RECT 293.460 295.700 295.540 296.660 ;
        RECT 0.700 4.300 295.540 295.700 ;
        RECT 1.140 3.500 12.860 4.300 ;
        RECT 14.580 3.500 26.300 4.300 ;
        RECT 28.020 3.500 43.100 4.300 ;
        RECT 44.820 3.500 56.540 4.300 ;
        RECT 58.260 3.500 73.340 4.300 ;
        RECT 75.060 3.500 86.780 4.300 ;
        RECT 88.500 3.500 103.580 4.300 ;
        RECT 105.300 3.500 117.020 4.300 ;
        RECT 118.740 3.500 133.820 4.300 ;
        RECT 135.540 3.500 147.260 4.300 ;
        RECT 148.980 3.500 160.700 4.300 ;
        RECT 162.420 3.500 177.500 4.300 ;
        RECT 179.220 3.500 190.940 4.300 ;
        RECT 192.660 3.500 207.740 4.300 ;
        RECT 209.460 3.500 221.180 4.300 ;
        RECT 222.900 3.500 237.980 4.300 ;
        RECT 239.700 3.500 251.420 4.300 ;
        RECT 253.140 3.500 268.220 4.300 ;
        RECT 269.940 3.500 281.660 4.300 ;
        RECT 283.380 3.500 295.100 4.300 ;
      LAYER Metal3 ;
        RECT 3.640 291.740 295.700 292.180 ;
        RECT 3.640 283.380 296.660 291.740 ;
        RECT 4.300 281.660 296.660 283.380 ;
        RECT 3.640 280.020 296.660 281.660 ;
        RECT 3.640 278.300 295.700 280.020 ;
        RECT 3.640 266.580 296.660 278.300 ;
        RECT 4.300 264.860 296.660 266.580 ;
        RECT 3.640 263.220 296.660 264.860 ;
        RECT 3.640 261.500 295.700 263.220 ;
        RECT 3.640 253.140 296.660 261.500 ;
        RECT 4.300 251.420 296.660 253.140 ;
        RECT 3.640 249.780 296.660 251.420 ;
        RECT 3.640 248.060 295.700 249.780 ;
        RECT 3.640 239.700 296.660 248.060 ;
        RECT 4.300 237.980 296.660 239.700 ;
        RECT 3.640 236.340 296.660 237.980 ;
        RECT 3.640 234.620 295.700 236.340 ;
        RECT 3.640 222.900 296.660 234.620 ;
        RECT 4.300 221.180 296.660 222.900 ;
        RECT 3.640 219.540 296.660 221.180 ;
        RECT 3.640 217.820 295.700 219.540 ;
        RECT 3.640 209.460 296.660 217.820 ;
        RECT 4.300 207.740 296.660 209.460 ;
        RECT 3.640 206.100 296.660 207.740 ;
        RECT 3.640 204.380 295.700 206.100 ;
        RECT 3.640 192.660 296.660 204.380 ;
        RECT 4.300 190.940 296.660 192.660 ;
        RECT 3.640 189.300 296.660 190.940 ;
        RECT 3.640 187.580 295.700 189.300 ;
        RECT 3.640 179.220 296.660 187.580 ;
        RECT 4.300 177.500 296.660 179.220 ;
        RECT 3.640 175.860 296.660 177.500 ;
        RECT 3.640 174.140 295.700 175.860 ;
        RECT 3.640 162.420 296.660 174.140 ;
        RECT 4.300 160.700 296.660 162.420 ;
        RECT 3.640 159.060 296.660 160.700 ;
        RECT 3.640 157.340 295.700 159.060 ;
        RECT 3.640 148.980 296.660 157.340 ;
        RECT 4.300 147.260 296.660 148.980 ;
        RECT 3.640 145.620 296.660 147.260 ;
        RECT 3.640 143.900 295.700 145.620 ;
        RECT 3.640 132.180 296.660 143.900 ;
        RECT 4.300 130.460 296.660 132.180 ;
        RECT 3.640 128.820 296.660 130.460 ;
        RECT 3.640 127.100 295.700 128.820 ;
        RECT 3.640 118.740 296.660 127.100 ;
        RECT 4.300 117.020 296.660 118.740 ;
        RECT 3.640 115.380 296.660 117.020 ;
        RECT 3.640 113.660 295.700 115.380 ;
        RECT 3.640 105.300 296.660 113.660 ;
        RECT 4.300 103.580 296.660 105.300 ;
        RECT 3.640 101.940 296.660 103.580 ;
        RECT 3.640 100.220 295.700 101.940 ;
        RECT 3.640 88.500 296.660 100.220 ;
        RECT 4.300 86.780 296.660 88.500 ;
        RECT 3.640 85.140 296.660 86.780 ;
        RECT 3.640 83.420 295.700 85.140 ;
        RECT 3.640 75.060 296.660 83.420 ;
        RECT 4.300 73.340 296.660 75.060 ;
        RECT 3.640 71.700 296.660 73.340 ;
        RECT 3.640 69.980 295.700 71.700 ;
        RECT 3.640 58.260 296.660 69.980 ;
        RECT 4.300 56.540 296.660 58.260 ;
        RECT 3.640 54.900 296.660 56.540 ;
        RECT 3.640 53.180 295.700 54.900 ;
        RECT 3.640 44.820 296.660 53.180 ;
        RECT 4.300 43.100 296.660 44.820 ;
        RECT 3.640 41.460 296.660 43.100 ;
        RECT 3.640 39.740 295.700 41.460 ;
        RECT 3.640 28.020 296.660 39.740 ;
        RECT 4.300 26.300 296.660 28.020 ;
        RECT 3.640 24.660 296.660 26.300 ;
        RECT 3.640 22.940 295.700 24.660 ;
        RECT 3.640 14.580 296.660 22.940 ;
        RECT 4.300 12.860 296.660 14.580 ;
        RECT 3.640 11.220 296.660 12.860 ;
        RECT 3.640 10.780 295.700 11.220 ;
      LAYER Metal4 ;
        RECT 24.220 118.250 98.740 231.750 ;
        RECT 100.940 118.250 175.540 231.750 ;
        RECT 177.740 118.250 197.540 231.750 ;
  END
END cntr_example
END LIBRARY

