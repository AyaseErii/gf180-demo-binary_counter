// This is the unpowered netlist.
module cntr_example (wb_clk_i,
    wb_rst_i,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire clknet_0_wb_clk_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _253_ (.A1(net52),
    .A2(net49),
    .A3(_100_),
    .A4(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _254_ (.A1(net63),
    .A2(net64),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _255_ (.A1(net66),
    .A2(net65),
    .A3(_065_),
    .A4(_103_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _256_ (.I(net43),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _257_ (.I(net40),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _258_ (.A1(net42),
    .A2(net41),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _259_ (.A1(net39),
    .A2(net38),
    .A3(net68),
    .A4(net67),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _260_ (.A1(_105_),
    .A2(_106_),
    .A3(_107_),
    .A4(_108_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _261_ (.A1(_102_),
    .A2(_104_),
    .A3(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _262_ (.A1(net58),
    .A2(net57),
    .A3(_099_),
    .A4(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _263_ (.I(net61),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _264_ (.A1(net60),
    .A2(_111_),
    .B(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _265_ (.A1(_112_),
    .A2(net60),
    .A3(_111_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _266_ (.A1(net36),
    .A2(_113_),
    .A3(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _267_ (.A1(_073_),
    .A2(net25),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _268_ (.A1(_071_),
    .A2(_115_),
    .A3(_116_),
    .B1(_112_),
    .B2(_082_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _269_ (.A1(net60),
    .A2(_111_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _270_ (.A1(_076_),
    .A2(_117_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _271_ (.A1(_073_),
    .A2(net24),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _272_ (.I(net60),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _273_ (.A1(_071_),
    .A2(_118_),
    .A3(_119_),
    .B1(_120_),
    .B2(_082_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _274_ (.I(net58),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _275_ (.A1(net57),
    .A2(_099_),
    .A3(_110_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _276_ (.A1(_121_),
    .A2(_122_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _277_ (.A1(_076_),
    .A2(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _278_ (.A1(_073_),
    .A2(net22),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _279_ (.A1(_071_),
    .A2(_124_),
    .A3(_125_),
    .B1(_121_),
    .B2(_082_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _280_ (.I(_070_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _281_ (.I(net57),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _282_ (.A1(_099_),
    .A2(_110_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _283_ (.A1(_127_),
    .A2(_128_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _284_ (.A1(_076_),
    .A2(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _285_ (.A1(_073_),
    .A2(net21),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _286_ (.A1(_126_),
    .A2(_130_),
    .A3(_131_),
    .B1(_127_),
    .B2(_082_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _287_ (.A1(net55),
    .A2(net54),
    .A3(net53),
    .A4(_110_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _288_ (.A1(net56),
    .A2(_132_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _289_ (.A1(_076_),
    .A2(_133_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _290_ (.A1(_073_),
    .A2(net20),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _291_ (.A1(_126_),
    .A2(_134_),
    .A3(_135_),
    .B1(_095_),
    .B2(_082_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _292_ (.A1(net52),
    .A2(net49),
    .A3(_100_),
    .A4(_101_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _293_ (.A1(net66),
    .A2(net65),
    .A3(_065_),
    .A4(_103_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _294_ (.I(net39),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _295_ (.I(net38),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _296_ (.A1(net43),
    .A2(net40),
    .A3(net68),
    .A4(net67),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _297_ (.A1(_138_),
    .A2(_139_),
    .A3(_107_),
    .A4(_140_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _298_ (.A1(net53),
    .A2(_136_),
    .A3(_137_),
    .A4(_141_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _299_ (.A1(net54),
    .A2(_142_),
    .B(net55),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _300_ (.A1(_132_),
    .A2(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _301_ (.A1(_076_),
    .A2(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _302_ (.I(_072_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _303_ (.A1(_146_),
    .A2(net19),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _304_ (.A1(_126_),
    .A2(_145_),
    .A3(_147_),
    .B1(_096_),
    .B2(_082_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _305_ (.A1(_097_),
    .A2(_142_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _306_ (.A1(_072_),
    .A2(_148_),
    .Z(_149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _307_ (.A1(_146_),
    .A2(net18),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _308_ (.I(_068_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _309_ (.A1(_126_),
    .A2(_149_),
    .A3(_150_),
    .B1(_097_),
    .B2(_151_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _310_ (.A1(net53),
    .A2(_110_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _311_ (.A1(_076_),
    .A2(_152_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _312_ (.A1(_146_),
    .A2(net17),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _313_ (.A1(_126_),
    .A2(_153_),
    .A3(_154_),
    .B1(_098_),
    .B2(_151_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _314_ (.I(net52),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _315_ (.A1(net49),
    .A2(_101_),
    .A3(_137_),
    .A4(_141_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _316_ (.A1(net51),
    .A2(net50),
    .A3(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _317_ (.A1(_155_),
    .A2(_157_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _318_ (.A1(_064_),
    .A2(_158_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _319_ (.A1(_146_),
    .A2(net16),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _320_ (.A1(_126_),
    .A2(_159_),
    .A3(_160_),
    .B1(_155_),
    .B2(_151_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _321_ (.I(net51),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _322_ (.A1(net50),
    .A2(_156_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _323_ (.A1(_161_),
    .A2(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _324_ (.A1(_064_),
    .A2(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _325_ (.A1(_146_),
    .A2(net15),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _326_ (.A1(_126_),
    .A2(_164_),
    .A3(_165_),
    .B1(_161_),
    .B2(_151_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _327_ (.A1(net50),
    .A2(_156_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _328_ (.A1(_162_),
    .A2(_166_),
    .B(_064_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _329_ (.A1(_146_),
    .A2(net14),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _330_ (.I(net50),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _331_ (.A1(_126_),
    .A2(_167_),
    .A3(_168_),
    .B1(_169_),
    .B2(_151_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _332_ (.I(net44),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _333_ (.A1(net47),
    .A2(net46),
    .A3(net45),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _334_ (.A1(_170_),
    .A2(_171_),
    .A3(_104_),
    .A4(_109_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _335_ (.A1(net49),
    .A2(_172_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _336_ (.A1(_064_),
    .A2(_173_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _337_ (.A1(_146_),
    .A2(net13),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _338_ (.I(net49),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _339_ (.A1(_126_),
    .A2(_174_),
    .A3(_175_),
    .B1(_176_),
    .B2(_151_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _340_ (.I(_068_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _341_ (.I(net47),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _342_ (.A1(_104_),
    .A2(_109_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _343_ (.A1(net46),
    .A2(net45),
    .A3(net44),
    .A4(_179_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _344_ (.A1(_178_),
    .A2(_180_),
    .B(_172_),
    .C(net36),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _345_ (.A1(_076_),
    .A2(net11),
    .B(_181_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _346_ (.A1(_177_),
    .A2(_178_),
    .B1(_071_),
    .B2(_182_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _347_ (.I(net46),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _348_ (.A1(net45),
    .A2(net44),
    .A3(_179_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _349_ (.A1(_183_),
    .A2(_184_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _350_ (.A1(_180_),
    .A2(_185_),
    .B(_064_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _351_ (.A1(_146_),
    .A2(net10),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _352_ (.A1(_126_),
    .A2(_186_),
    .A3(_187_),
    .B1(_183_),
    .B2(_151_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _353_ (.I(_070_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _354_ (.I(net45),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _355_ (.A1(net44),
    .A2(_179_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _356_ (.A1(_189_),
    .A2(_190_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _357_ (.I(net36),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _358_ (.A1(_184_),
    .A2(_191_),
    .B(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _359_ (.A1(_146_),
    .A2(net9),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _360_ (.A1(_188_),
    .A2(_193_),
    .A3(_194_),
    .B1(_189_),
    .B2(_151_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _361_ (.A1(_104_),
    .A2(_109_),
    .B(_170_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _362_ (.A1(_190_),
    .A2(_195_),
    .B(_192_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _363_ (.A1(_146_),
    .A2(net8),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _364_ (.A1(_188_),
    .A2(_196_),
    .A3(_197_),
    .B1(_170_),
    .B2(_151_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _365_ (.A1(_104_),
    .A2(_108_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _366_ (.A1(net42),
    .A2(net41),
    .A3(net40),
    .A4(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _367_ (.A1(_105_),
    .A2(_199_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _368_ (.A1(_064_),
    .A2(_200_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _369_ (.I(_072_),
    .Z(_202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _370_ (.A1(_202_),
    .A2(net7),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _371_ (.A1(_188_),
    .A2(_201_),
    .A3(_203_),
    .B1(_105_),
    .B2(_151_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _372_ (.I(net42),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _373_ (.A1(net41),
    .A2(net40),
    .A3(_198_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _374_ (.A1(_204_),
    .A2(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _375_ (.A1(_199_),
    .A2(_206_),
    .B(_192_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _376_ (.A1(_202_),
    .A2(net6),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _377_ (.A1(_188_),
    .A2(_207_),
    .A3(_208_),
    .B1(_204_),
    .B2(_177_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _378_ (.I(net41),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _379_ (.A1(net40),
    .A2(_198_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _380_ (.A1(_209_),
    .A2(_210_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _381_ (.A1(_205_),
    .A2(_211_),
    .B(_192_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _382_ (.A1(_202_),
    .A2(net5),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _383_ (.A1(_188_),
    .A2(_212_),
    .A3(_213_),
    .B1(_209_),
    .B2(_177_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _384_ (.A1(_104_),
    .A2(_108_),
    .B(_106_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _385_ (.A1(_210_),
    .A2(_214_),
    .B(_192_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _386_ (.A1(_202_),
    .A2(net4),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _387_ (.A1(_188_),
    .A2(_215_),
    .A3(_216_),
    .B1(_106_),
    .B2(_177_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _388_ (.A1(net68),
    .A2(net67),
    .A3(_137_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _389_ (.A1(_139_),
    .A2(_217_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _390_ (.A1(_138_),
    .A2(_218_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _391_ (.A1(_064_),
    .A2(_219_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _392_ (.A1(_202_),
    .A2(net3),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _393_ (.A1(_188_),
    .A2(_220_),
    .A3(_221_),
    .B1(_138_),
    .B2(_177_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _394_ (.A1(_139_),
    .A2(_217_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _395_ (.A1(_218_),
    .A2(_222_),
    .B(_192_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _396_ (.A1(_202_),
    .A2(net2),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _397_ (.A1(_188_),
    .A2(_223_),
    .A3(_224_),
    .B1(_139_),
    .B2(_177_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _398_ (.I(net68),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _399_ (.A1(net67),
    .A2(_137_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _400_ (.A1(_225_),
    .A2(_226_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _401_ (.A1(_217_),
    .A2(_227_),
    .B(_192_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _402_ (.A1(_202_),
    .A2(net32),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _403_ (.A1(_188_),
    .A2(_228_),
    .A3(_229_),
    .B1(_225_),
    .B2(_177_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _404_ (.I(net67),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _405_ (.A1(_230_),
    .A2(_104_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _406_ (.A1(_226_),
    .A2(_231_),
    .B(_192_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _407_ (.A1(_202_),
    .A2(net31),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _408_ (.A1(_188_),
    .A2(_232_),
    .A3(_233_),
    .B1(_230_),
    .B2(_177_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _409_ (.I(net66),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _410_ (.A1(net65),
    .A2(_065_),
    .A3(_103_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _411_ (.A1(_234_),
    .A2(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _412_ (.A1(_072_),
    .A2(_104_),
    .A3(_236_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _413_ (.A1(_076_),
    .A2(net30),
    .B(_237_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _414_ (.A1(_068_),
    .A2(_234_),
    .B1(_071_),
    .B2(_238_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _415_ (.I(net65),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _416_ (.A1(_065_),
    .A2(_103_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _417_ (.A1(_239_),
    .A2(_240_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _418_ (.A1(_235_),
    .A2(_241_),
    .B(_192_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _419_ (.A1(_202_),
    .A2(net29),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _420_ (.A1(_070_),
    .A2(_242_),
    .A3(_243_),
    .B1(_239_),
    .B2(_177_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _421_ (.A1(net63),
    .A2(_065_),
    .B(net64),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _422_ (.I(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _423_ (.A1(_240_),
    .A2(_245_),
    .B(_192_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _424_ (.A1(_202_),
    .A2(net28),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _425_ (.I(net64),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _426_ (.A1(_070_),
    .A2(_246_),
    .A3(_247_),
    .B1(_248_),
    .B2(_177_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _427_ (.I(net33),
    .Z(_249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _428_ (.I(_249_),
    .Z(_250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _429_ (.I(_250_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _430_ (.I(_250_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _431_ (.I(_250_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _432_ (.I(_250_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _433_ (.I(_250_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _434_ (.I(_250_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _435_ (.I(_250_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _436_ (.I(_250_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _437_ (.I(_250_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _438_ (.I(_250_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _439_ (.I(_249_),
    .Z(_251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _440_ (.I(_251_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _441_ (.I(_251_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _442_ (.I(_251_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _443_ (.I(_251_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _444_ (.I(_251_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _445_ (.I(_251_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _446_ (.I(_251_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _447_ (.I(_251_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _448_ (.I(_251_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _449_ (.I(_251_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _450_ (.I(_249_),
    .Z(_252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _451_ (.I(_252_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _452_ (.I(_252_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _453_ (.I(_252_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _454_ (.I(_252_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _455_ (.I(_252_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _456_ (.I(_252_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _457_ (.I(_252_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _458_ (.I(_252_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _459_ (.I(_252_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _460_ (.I(_252_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _461_ (.I(_249_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _462_ (.I(_249_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _463_ (.I(net36),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _464_ (.A1(net62),
    .A2(net59),
    .A3(net48),
    .A4(net37),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _465_ (.A1(net63),
    .A2(_065_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _466_ (.A1(_064_),
    .A2(_066_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _467_ (.I(net34),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _468_ (.I(net35),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _469_ (.A1(_068_),
    .A2(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _470_ (.I(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _471_ (.I(net36),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _472_ (.I(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _473_ (.A1(_073_),
    .A2(net27),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _474_ (.I(net63),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _475_ (.A1(_067_),
    .A2(_071_),
    .A3(_074_),
    .B1(_068_),
    .B2(_075_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _476_ (.I(net36),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _477_ (.I(net62),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _478_ (.A1(net59),
    .A2(net48),
    .A3(net37),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _479_ (.A1(_077_),
    .A2(_078_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _480_ (.A1(_076_),
    .A2(_079_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _481_ (.A1(_073_),
    .A2(net26),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _482_ (.I(_068_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _483_ (.A1(_071_),
    .A2(_080_),
    .A3(_081_),
    .B1(_077_),
    .B2(_082_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _484_ (.I(net59),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _485_ (.A1(net48),
    .A2(net37),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _486_ (.A1(_083_),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _487_ (.A1(_078_),
    .A2(_085_),
    .B(_064_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _488_ (.A1(_073_),
    .A2(net23),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _489_ (.A1(_071_),
    .A2(_086_),
    .A3(_087_),
    .B1(_083_),
    .B2(_082_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _490_ (.I(net48),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _491_ (.I(net37),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _492_ (.A1(_088_),
    .A2(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _493_ (.A1(_084_),
    .A2(_090_),
    .B(_064_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _494_ (.A1(_073_),
    .A2(net12),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _495_ (.A1(_071_),
    .A2(_091_),
    .A3(_092_),
    .B1(_088_),
    .B2(_082_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _496_ (.A1(_089_),
    .A2(_076_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _497_ (.A1(net1),
    .A2(_073_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _498_ (.A1(_071_),
    .A2(_093_),
    .A3(_094_),
    .B1(_089_),
    .B2(_082_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _499_ (.I(net56),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _500_ (.I(net55),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _501_ (.I(net54),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _502_ (.I(net53),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _503_ (.A1(_095_),
    .A2(_096_),
    .A3(_097_),
    .A4(_098_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _504_ (.A1(net51),
    .A2(net50),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _505_ (.A1(net47),
    .A2(net46),
    .A3(net45),
    .A4(net44),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _506_ (.D(_032_),
    .RN(_000_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _507_ (.D(_033_),
    .RN(_001_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _508_ (.D(_034_),
    .RN(_002_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _509_ (.D(_035_),
    .RN(_003_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _510_ (.D(_036_),
    .RN(_004_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _511_ (.D(_037_),
    .RN(_005_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _512_ (.D(_038_),
    .RN(_006_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _513_ (.D(_039_),
    .RN(_007_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _514_ (.D(_040_),
    .RN(_008_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _515_ (.D(_041_),
    .RN(_009_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _516_ (.D(_042_),
    .RN(_010_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _517_ (.D(_043_),
    .RN(_011_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _518_ (.D(_044_),
    .RN(_012_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _519_ (.D(_045_),
    .RN(_013_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _520_ (.D(_046_),
    .RN(_014_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _521_ (.D(_047_),
    .RN(_015_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _522_ (.D(_048_),
    .RN(_016_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _523_ (.D(_049_),
    .RN(_017_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _524_ (.D(_050_),
    .RN(_018_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _525_ (.D(_051_),
    .RN(_019_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _526_ (.D(_052_),
    .RN(_020_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _527_ (.D(_053_),
    .RN(_021_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _528_ (.D(_054_),
    .RN(_022_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _529_ (.D(_055_),
    .RN(_023_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _530_ (.D(_056_),
    .RN(_024_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _531_ (.D(_057_),
    .RN(_025_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _532_ (.D(_058_),
    .RN(_026_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _533_ (.D(_059_),
    .RN(_027_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _534_ (.D(_060_),
    .RN(_028_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _535_ (.D(_061_),
    .RN(_029_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _536_ (.D(_062_),
    .RN(_030_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _537_ (.D(_063_),
    .RN(_031_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(io_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(io_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(io_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(io_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(io_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(io_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(io_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(io_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(io_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(io_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(io_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(io_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(io_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(io_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(io_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(io_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(io_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(io_in[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(io_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(io_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(io_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(io_in[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(io_in[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(io_in[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(wb_rst_i),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(wbs_cyc_i),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(wbs_stb_i),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(wbs_we_i),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output38 (.I(net38),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output39 (.I(net39),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output40 (.I(net40),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output42 (.I(net42),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output50 (.I(net50),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output52 (.I(net52),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output53 (.I(net53),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output54 (.I(net54),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output55 (.I(net55),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output56 (.I(net56),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output58 (.I(net58),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output59 (.I(net59),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output65 (.I(net65),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output67 (.I(net67),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output68 (.I(net68),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__RN (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__RN (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__RN (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__RN (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__RN (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__RN (.I(_008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__RN (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__RN (.I(_010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__RN (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__RN (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__RN (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__RN (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__RN (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__RN (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__RN (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__RN (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__RN (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__RN (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__RN (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__RN (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__RN (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__RN (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__RN (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__RN (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__RN (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__RN (.I(_031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__D (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__D (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__D (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__D (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__D (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__D (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__D (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__D (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__D (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__D (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__D (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__D (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__D (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__D (.I(_045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__D (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__D (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__D (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__D (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__D (.I(_050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__D (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__D (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__D (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__D (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__D (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__D (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__D (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__D (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__D (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__D (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__D (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__D (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__D (.I(_063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__B (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__B (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__B (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__B (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A3 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A3 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A1 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__I (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__B1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__I (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__I (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__I (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__I (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A2 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__B1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__B1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A3 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__B2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A3 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A3 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__B1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A2 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__B1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A3 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__B1 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A1 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A4 (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__B1 (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A1 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A2 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A3 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__A1 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A3 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__B1 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__A1 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A1 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A3 (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A3 (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A2 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__A2 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A4 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A2 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__A2 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A4 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A3 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__A2 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A4 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A2 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A3 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A4 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A2 (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A3 (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A2 (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__B1 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A1 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__B (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A2 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__A2 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A1 (.I(_132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__A2 (.I(_132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A2 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A2 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A3 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A3 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A3 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__B1 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__A1 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A1 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__B1 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A1 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A1 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A4 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A4 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A2 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A2 (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A1 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A3 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__A2 (.I(_149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__B2 (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__A3 (.I(_154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A2 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A2 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A3 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A3 (.I(_160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__A3 (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A3 (.I(_168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__B1 (.I(_170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__B (.I(_170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A1 (.I(_170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__B (.I(_172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A2 (.I(_172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__B2 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A1 (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__A1 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__A2 (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__B1 (.I(_183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__A1 (.I(_183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__A1 (.I(_184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__A2 (.I(_184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__A1 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__A2 (.I(_190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__B (.I(_192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__A3 (.I(_194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A3 (.I(_197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__A1 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__A2 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A1 (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__A3 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__B1 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__A1 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__A3 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A3 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A2 (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A1 (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__A1 (.I(_235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A2 (.I(_235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A3 (.I(_236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__B2 (.I(_238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A1 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__A2 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A3 (.I(_243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__I (.I(_249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(_249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__I (.I(_249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__I (.I(_249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__I (.I(_249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__431__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__I (.I(_250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__I (.I(_251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__I (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(io_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__C (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__A3 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A4 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A3 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A4 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__A2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A3 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A3 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A3 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A3 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A3 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__B (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__B (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A2 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A2 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A4 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__A4 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A3 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__A3 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__CLK (.I(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__CLK (.I(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_508 ();
 assign io_out[32] = net69;
 assign io_out[33] = net70;
 assign io_out[34] = net71;
 assign io_out[35] = net72;
 assign io_out[36] = net73;
 assign io_out[37] = net74;
endmodule

